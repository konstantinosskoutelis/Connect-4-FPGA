module winner_sprite(
  input logic[12:0] addr,
	output logic data
);

logic[4859:0] mem;

//Custom Memory For Winner Sprite
always_comb begin
mem[0] = 0;
mem[1] = 0;
mem[2] = 0;
mem[3] = 0;
mem[4] = 0;
mem[5] = 0;
mem[6] = 0;
mem[7] = 0;
mem[8] = 0;
mem[9] = 0;
mem[10] = 0;
mem[11] = 0;
mem[12] = 0;
mem[13] = 0;
mem[14] = 0;
mem[15] = 0;
mem[16] = 0;
mem[17] = 0;
mem[18] = 0;
mem[19] = 0;
mem[20] = 0;
mem[21] = 1;
mem[22] = 1;
mem[23] = 1;
mem[24] = 0;
mem[25] = 0;
mem[26] = 0;
mem[27] = 0;
mem[28] = 0;
mem[29] = 0;
mem[30] = 0;
mem[31] = 0;
mem[32] = 0;
mem[33] = 0;
mem[34] = 1;
mem[35] = 1;
mem[36] = 0;
mem[37] = 0;
mem[38] = 0;
mem[39] = 0;
mem[40] = 0;
mem[41] = 0;
mem[42] = 0;
mem[43] = 0;
mem[44] = 0;
mem[45] = 0;
mem[46] = 1;
mem[47] = 1;
mem[48] = 1;
mem[49] = 1;
mem[50] = 0;
mem[51] = 0;
mem[52] = 0;
mem[53] = 0;
mem[54] = 0;
mem[55] = 0;
mem[56] = 1;
mem[57] = 1;
mem[58] = 1;
mem[59] = 0;
mem[60] = 0;
mem[61] = 0;
mem[62] = 0;
mem[63] = 0;
mem[64] = 0;
mem[65] = 0;
mem[66] = 0;
mem[67] = 0;
mem[68] = 0;
mem[69] = 1;
mem[70] = 0;
mem[71] = 0;
mem[72] = 0;
mem[73] = 0;
mem[74] = 0;
mem[75] = 0;
mem[76] = 0;
mem[77] = 0;
mem[78] = 0;
mem[79] = 0;
mem[80] = 0;
mem[81] = 0;
mem[82] = 0;
mem[83] = 0;
mem[84] = 0;
mem[85] = 0;
mem[86] = 0;
mem[87] = 0;
mem[88] = 0;
mem[89] = 0;
mem[90] = 0;
mem[91] = 0;
mem[92] = 0;
mem[93] = 0;
mem[94] = 0;
mem[95] = 0;
mem[96] = 0;
mem[97] = 0;
mem[98] = 1;
mem[99] = 1;
mem[100] = 1;
mem[101] = 1;
mem[102] = 0;
mem[103] = 0;
mem[104] = 0;
mem[105] = 0;
mem[106] = 0;
mem[107] = 0;
mem[108] = 0;
mem[109] = 0;
mem[110] = 1;
mem[111] = 1;
mem[112] = 1;
mem[113] = 1;
mem[114] = 1;
mem[115] = 0;
mem[116] = 0;
mem[117] = 0;
mem[118] = 0;
mem[119] = 0;
mem[120] = 0;
mem[121] = 0;
mem[122] = 0;
mem[123] = 1;
mem[124] = 1;
mem[125] = 1;
mem[126] = 1;
mem[127] = 0;
mem[128] = 0;
mem[129] = 0;
mem[130] = 0;
mem[131] = 0;
mem[132] = 0;
mem[133] = 0;
mem[134] = 0;
mem[135] = 0;
mem[136] = 1;
mem[137] = 1;
mem[138] = 1;
mem[139] = 1;
mem[140] = 0;
mem[141] = 0;
mem[142] = 0;
mem[143] = 0;
mem[144] = 0;
mem[145] = 0;
mem[146] = 1;
mem[147] = 1;
mem[148] = 1;
mem[149] = 0;
mem[150] = 0;
mem[151] = 0;
mem[152] = 0;
mem[153] = 0;
mem[154] = 0;
mem[155] = 0;
mem[156] = 0;
mem[157] = 1;
mem[158] = 1;
mem[159] = 1;
mem[160] = 0;
mem[161] = 0;
mem[162] = 0;
mem[163] = 0;
mem[164] = 0;
mem[165] = 0;
mem[166] = 0;
mem[167] = 0;
mem[168] = 0;
mem[169] = 0;
mem[170] = 0;
mem[171] = 0;
mem[172] = 0;
mem[173] = 0;
mem[174] = 0;
mem[175] = 0;
mem[176] = 0;
mem[177] = 0;
mem[178] = 0;
mem[179] = 0;
mem[180] = 0;
mem[181] = 0;
mem[182] = 0;
mem[183] = 0;
mem[184] = 0;
mem[185] = 0;
mem[186] = 0;
mem[187] = 0;
mem[188] = 1;
mem[189] = 1;
mem[190] = 1;
mem[191] = 1;
mem[192] = 1;
mem[193] = 1;
mem[194] = 0;
mem[195] = 0;
mem[196] = 0;
mem[197] = 0;
mem[198] = 0;
mem[199] = 0;
mem[200] = 1;
mem[201] = 1;
mem[202] = 1;
mem[203] = 1;
mem[204] = 1;
mem[205] = 0;
mem[206] = 0;
mem[207] = 0;
mem[208] = 0;
mem[209] = 0;
mem[210] = 0;
mem[211] = 0;
mem[212] = 0;
mem[213] = 1;
mem[214] = 1;
mem[215] = 1;
mem[216] = 1;
mem[217] = 0;
mem[218] = 0;
mem[219] = 0;
mem[220] = 0;
mem[221] = 0;
mem[222] = 0;
mem[223] = 0;
mem[224] = 0;
mem[225] = 1;
mem[226] = 1;
mem[227] = 1;
mem[228] = 1;
mem[229] = 1;
mem[230] = 1;
mem[231] = 0;
mem[232] = 0;
mem[233] = 0;
mem[234] = 0;
mem[235] = 0;
mem[236] = 1;
mem[237] = 1;
mem[238] = 1;
mem[239] = 1;
mem[240] = 0;
mem[241] = 0;
mem[242] = 0;
mem[243] = 0;
mem[244] = 0;
mem[245] = 0;
mem[246] = 1;
mem[247] = 1;
mem[248] = 1;
mem[249] = 1;
mem[250] = 0;
mem[251] = 0;
mem[252] = 0;
mem[253] = 0;
mem[254] = 0;
mem[255] = 0;
mem[256] = 0;
mem[257] = 0;
mem[258] = 0;
mem[259] = 0;
mem[260] = 0;
mem[261] = 0;
mem[262] = 0;
mem[263] = 0;
mem[264] = 0;
mem[265] = 0;
mem[266] = 0;
mem[267] = 0;
mem[268] = 0;
mem[269] = 0;
mem[270] = 0;
mem[271] = 0;
mem[272] = 0;
mem[273] = 0;
mem[274] = 0;
mem[275] = 0;
mem[276] = 0;
mem[277] = 0;
mem[278] = 0;
mem[279] = 1;
mem[280] = 1;
mem[281] = 1;
mem[282] = 1;
mem[283] = 1;
mem[284] = 1;
mem[285] = 0;
mem[286] = 0;
mem[287] = 0;
mem[288] = 0;
mem[289] = 0;
mem[290] = 1;
mem[291] = 1;
mem[292] = 0;
mem[293] = 1;
mem[294] = 1;
mem[295] = 1;
mem[296] = 0;
mem[297] = 0;
mem[298] = 0;
mem[299] = 0;
mem[300] = 0;
mem[301] = 0;
mem[302] = 1;
mem[303] = 1;
mem[304] = 1;
mem[305] = 0;
mem[306] = 1;
mem[307] = 1;
mem[308] = 0;
mem[309] = 0;
mem[310] = 0;
mem[311] = 0;
mem[312] = 0;
mem[313] = 0;
mem[314] = 1;
mem[315] = 1;
mem[316] = 1;
mem[317] = 0;
mem[318] = 1;
mem[319] = 1;
mem[320] = 1;
mem[321] = 0;
mem[322] = 0;
mem[323] = 0;
mem[324] = 0;
mem[325] = 1;
mem[326] = 1;
mem[327] = 1;
mem[328] = 1;
mem[329] = 1;
mem[330] = 0;
mem[331] = 0;
mem[332] = 0;
mem[333] = 0;
mem[334] = 0;
mem[335] = 0;
mem[336] = 1;
mem[337] = 1;
mem[338] = 1;
mem[339] = 1;
mem[340] = 1;
mem[341] = 0;
mem[342] = 0;
mem[343] = 0;
mem[344] = 0;
mem[345] = 0;
mem[346] = 0;
mem[347] = 0;
mem[348] = 0;
mem[349] = 0;
mem[350] = 0;
mem[351] = 0;
mem[352] = 0;
mem[353] = 0;
mem[354] = 0;
mem[355] = 0;
mem[356] = 0;
mem[357] = 0;
mem[358] = 0;
mem[359] = 0;
mem[360] = 0;
mem[361] = 0;
mem[362] = 0;
mem[363] = 0;
mem[364] = 0;
mem[365] = 0;
mem[366] = 0;
mem[367] = 0;
mem[368] = 0;
mem[369] = 1;
mem[370] = 1;
mem[371] = 1;
mem[372] = 1;
mem[373] = 1;
mem[374] = 1;
mem[375] = 1;
mem[376] = 1;
mem[377] = 0;
mem[378] = 0;
mem[379] = 1;
mem[380] = 1;
mem[381] = 1;
mem[382] = 0;
mem[383] = 1;
mem[384] = 1;
mem[385] = 1;
mem[386] = 1;
mem[387] = 0;
mem[388] = 0;
mem[389] = 0;
mem[390] = 0;
mem[391] = 0;
mem[392] = 1;
mem[393] = 1;
mem[394] = 0;
mem[395] = 0;
mem[396] = 1;
mem[397] = 1;
mem[398] = 0;
mem[399] = 0;
mem[400] = 0;
mem[401] = 0;
mem[402] = 0;
mem[403] = 1;
mem[404] = 1;
mem[405] = 1;
mem[406] = 0;
mem[407] = 0;
mem[408] = 0;
mem[409] = 1;
mem[410] = 1;
mem[411] = 1;
mem[412] = 0;
mem[413] = 0;
mem[414] = 1;
mem[415] = 1;
mem[416] = 1;
mem[417] = 0;
mem[418] = 1;
mem[419] = 1;
mem[420] = 1;
mem[421] = 0;
mem[422] = 0;
mem[423] = 0;
mem[424] = 0;
mem[425] = 1;
mem[426] = 1;
mem[427] = 1;
mem[428] = 0;
mem[429] = 1;
mem[430] = 1;
mem[431] = 0;
mem[432] = 0;
mem[433] = 0;
mem[434] = 0;
mem[435] = 0;
mem[436] = 0;
mem[437] = 0;
mem[438] = 0;
mem[439] = 0;
mem[440] = 0;
mem[441] = 1;
mem[442] = 1;
mem[443] = 1;
mem[444] = 0;
mem[445] = 0;
mem[446] = 0;
mem[447] = 0;
mem[448] = 0;
mem[449] = 0;
mem[450] = 0;
mem[451] = 0;
mem[452] = 0;
mem[453] = 0;
mem[454] = 0;
mem[455] = 0;
mem[456] = 0;
mem[457] = 0;
mem[458] = 0;
mem[459] = 0;
mem[460] = 1;
mem[461] = 1;
mem[462] = 0;
mem[463] = 0;
mem[464] = 1;
mem[465] = 1;
mem[466] = 1;
mem[467] = 1;
mem[468] = 1;
mem[469] = 1;
mem[470] = 1;
mem[471] = 0;
mem[472] = 0;
mem[473] = 0;
mem[474] = 1;
mem[475] = 1;
mem[476] = 1;
mem[477] = 0;
mem[478] = 0;
mem[479] = 0;
mem[480] = 0;
mem[481] = 1;
mem[482] = 1;
mem[483] = 1;
mem[484] = 0;
mem[485] = 0;
mem[486] = 0;
mem[487] = 1;
mem[488] = 1;
mem[489] = 0;
mem[490] = 0;
mem[491] = 0;
mem[492] = 0;
mem[493] = 1;
mem[494] = 1;
mem[495] = 0;
mem[496] = 0;
mem[497] = 0;
mem[498] = 0;
mem[499] = 0;
mem[500] = 1;
mem[501] = 1;
mem[502] = 0;
mem[503] = 1;
mem[504] = 1;
mem[505] = 1;
mem[506] = 0;
mem[507] = 0;
mem[508] = 1;
mem[509] = 1;
mem[510] = 1;
mem[511] = 0;
mem[512] = 0;
mem[513] = 0;
mem[514] = 1;
mem[515] = 1;
mem[516] = 1;
mem[517] = 0;
mem[518] = 0;
mem[519] = 1;
mem[520] = 1;
mem[521] = 0;
mem[522] = 0;
mem[523] = 0;
mem[524] = 0;
mem[525] = 0;
mem[526] = 0;
mem[527] = 0;
mem[528] = 0;
mem[529] = 1;
mem[530] = 1;
mem[531] = 1;
mem[532] = 1;
mem[533] = 1;
mem[534] = 1;
mem[535] = 0;
mem[536] = 0;
mem[537] = 0;
mem[538] = 0;
mem[539] = 0;
mem[540] = 0;
mem[541] = 0;
mem[542] = 0;
mem[543] = 0;
mem[544] = 0;
mem[545] = 0;
mem[546] = 0;
mem[547] = 0;
mem[548] = 0;
mem[549] = 0;
mem[550] = 1;
mem[551] = 1;
mem[552] = 1;
mem[553] = 0;
mem[554] = 0;
mem[555] = 0;
mem[556] = 1;
mem[557] = 1;
mem[558] = 1;
mem[559] = 1;
mem[560] = 1;
mem[561] = 0;
mem[562] = 0;
mem[563] = 0;
mem[564] = 1;
mem[565] = 1;
mem[566] = 1;
mem[567] = 0;
mem[568] = 0;
mem[569] = 0;
mem[570] = 0;
mem[571] = 1;
mem[572] = 1;
mem[573] = 0;
mem[574] = 0;
mem[575] = 0;
mem[576] = 0;
mem[577] = 1;
mem[578] = 1;
mem[579] = 0;
mem[580] = 0;
mem[581] = 0;
mem[582] = 1;
mem[583] = 1;
mem[584] = 1;
mem[585] = 0;
mem[586] = 0;
mem[587] = 0;
mem[588] = 0;
mem[589] = 0;
mem[590] = 1;
mem[591] = 1;
mem[592] = 1;
mem[593] = 1;
mem[594] = 0;
mem[595] = 0;
mem[596] = 0;
mem[597] = 0;
mem[598] = 1;
mem[599] = 1;
mem[600] = 1;
mem[601] = 0;
mem[602] = 0;
mem[603] = 0;
mem[604] = 1;
mem[605] = 1;
mem[606] = 1;
mem[607] = 0;
mem[608] = 0;
mem[609] = 1;
mem[610] = 1;
mem[611] = 1;
mem[612] = 0;
mem[613] = 0;
mem[614] = 0;
mem[615] = 0;
mem[616] = 0;
mem[617] = 0;
mem[618] = 1;
mem[619] = 1;
mem[620] = 1;
mem[621] = 1;
mem[622] = 1;
mem[623] = 1;
mem[624] = 0;
mem[625] = 0;
mem[626] = 0;
mem[627] = 0;
mem[628] = 0;
mem[629] = 0;
mem[630] = 0;
mem[631] = 0;
mem[632] = 0;
mem[633] = 0;
mem[634] = 0;
mem[635] = 0;
mem[636] = 0;
mem[637] = 0;
mem[638] = 0;
mem[639] = 0;
mem[640] = 1;
mem[641] = 1;
mem[642] = 1;
mem[643] = 0;
mem[644] = 0;
mem[645] = 0;
mem[646] = 0;
mem[647] = 1;
mem[648] = 1;
mem[649] = 1;
mem[650] = 0;
mem[651] = 0;
mem[652] = 0;
mem[653] = 0;
mem[654] = 1;
mem[655] = 1;
mem[656] = 1;
mem[657] = 0;
mem[658] = 0;
mem[659] = 0;
mem[660] = 1;
mem[661] = 1;
mem[662] = 1;
mem[663] = 0;
mem[664] = 0;
mem[665] = 0;
mem[666] = 0;
mem[667] = 0;
mem[668] = 1;
mem[669] = 1;
mem[670] = 0;
mem[671] = 1;
mem[672] = 1;
mem[673] = 1;
mem[674] = 0;
mem[675] = 0;
mem[676] = 0;
mem[677] = 0;
mem[678] = 0;
mem[679] = 0;
mem[680] = 0;
mem[681] = 1;
mem[682] = 1;
mem[683] = 1;
mem[684] = 1;
mem[685] = 0;
mem[686] = 0;
mem[687] = 0;
mem[688] = 0;
mem[689] = 1;
mem[690] = 1;
mem[691] = 1;
mem[692] = 0;
mem[693] = 1;
mem[694] = 1;
mem[695] = 1;
mem[696] = 0;
mem[697] = 0;
mem[698] = 0;
mem[699] = 0;
mem[700] = 1;
mem[701] = 1;
mem[702] = 0;
mem[703] = 0;
mem[704] = 0;
mem[705] = 0;
mem[706] = 0;
mem[707] = 1;
mem[708] = 1;
mem[709] = 1;
mem[710] = 0;
mem[711] = 1;
mem[712] = 1;
mem[713] = 0;
mem[714] = 0;
mem[715] = 0;
mem[716] = 0;
mem[717] = 0;
mem[718] = 0;
mem[719] = 0;
mem[720] = 0;
mem[721] = 0;
mem[722] = 0;
mem[723] = 0;
mem[724] = 0;
mem[725] = 0;
mem[726] = 0;
mem[727] = 0;
mem[728] = 0;
mem[729] = 0;
mem[730] = 1;
mem[731] = 1;
mem[732] = 1;
mem[733] = 0;
mem[734] = 0;
mem[735] = 0;
mem[736] = 0;
mem[737] = 0;
mem[738] = 0;
mem[739] = 0;
mem[740] = 0;
mem[741] = 0;
mem[742] = 0;
mem[743] = 0;
mem[744] = 0;
mem[745] = 0;
mem[746] = 1;
mem[747] = 1;
mem[748] = 0;
mem[749] = 1;
mem[750] = 1;
mem[751] = 1;
mem[752] = 0;
mem[753] = 0;
mem[754] = 0;
mem[755] = 0;
mem[756] = 0;
mem[757] = 0;
mem[758] = 1;
mem[759] = 1;
mem[760] = 1;
mem[761] = 1;
mem[762] = 1;
mem[763] = 0;
mem[764] = 0;
mem[765] = 0;
mem[766] = 0;
mem[767] = 0;
mem[768] = 0;
mem[769] = 0;
mem[770] = 0;
mem[771] = 1;
mem[772] = 1;
mem[773] = 0;
mem[774] = 0;
mem[775] = 0;
mem[776] = 0;
mem[777] = 0;
mem[778] = 0;
mem[779] = 1;
mem[780] = 1;
mem[781] = 1;
mem[782] = 1;
mem[783] = 1;
mem[784] = 0;
mem[785] = 0;
mem[786] = 0;
mem[787] = 0;
mem[788] = 0;
mem[789] = 0;
mem[790] = 1;
mem[791] = 1;
mem[792] = 1;
mem[793] = 0;
mem[794] = 0;
mem[795] = 0;
mem[796] = 1;
mem[797] = 1;
mem[798] = 1;
mem[799] = 0;
mem[800] = 0;
mem[801] = 1;
mem[802] = 1;
mem[803] = 0;
mem[804] = 0;
mem[805] = 0;
mem[806] = 0;
mem[807] = 0;
mem[808] = 0;
mem[809] = 0;
mem[810] = 0;
mem[811] = 0;
mem[812] = 0;
mem[813] = 0;
mem[814] = 0;
mem[815] = 0;
mem[816] = 0;
mem[817] = 0;
mem[818] = 0;
mem[819] = 0;
mem[820] = 0;
mem[821] = 1;
mem[822] = 1;
mem[823] = 1;
mem[824] = 0;
mem[825] = 0;
mem[826] = 0;
mem[827] = 0;
mem[828] = 0;
mem[829] = 0;
mem[830] = 0;
mem[831] = 0;
mem[832] = 0;
mem[833] = 0;
mem[834] = 0;
mem[835] = 1;
mem[836] = 1;
mem[837] = 1;
mem[838] = 0;
mem[839] = 0;
mem[840] = 1;
mem[841] = 1;
mem[842] = 0;
mem[843] = 0;
mem[844] = 0;
mem[845] = 0;
mem[846] = 0;
mem[847] = 0;
mem[848] = 0;
mem[849] = 1;
mem[850] = 1;
mem[851] = 1;
mem[852] = 1;
mem[853] = 0;
mem[854] = 0;
mem[855] = 0;
mem[856] = 0;
mem[857] = 0;
mem[858] = 0;
mem[859] = 0;
mem[860] = 0;
mem[861] = 0;
mem[862] = 0;
mem[863] = 0;
mem[864] = 0;
mem[865] = 0;
mem[866] = 0;
mem[867] = 0;
mem[868] = 0;
mem[869] = 0;
mem[870] = 1;
mem[871] = 1;
mem[872] = 1;
mem[873] = 0;
mem[874] = 0;
mem[875] = 0;
mem[876] = 0;
mem[877] = 0;
mem[878] = 0;
mem[879] = 0;
mem[880] = 0;
mem[881] = 0;
mem[882] = 1;
mem[883] = 0;
mem[884] = 1;
mem[885] = 1;
mem[886] = 1;
mem[887] = 1;
mem[888] = 0;
mem[889] = 0;
mem[890] = 0;
mem[891] = 1;
mem[892] = 1;
mem[893] = 0;
mem[894] = 0;
mem[895] = 0;
mem[896] = 0;
mem[897] = 0;
mem[898] = 0;
mem[899] = 0;
mem[900] = 0;
mem[901] = 0;
mem[902] = 0;
mem[903] = 0;
mem[904] = 0;
mem[905] = 0;
mem[906] = 0;
mem[907] = 0;
mem[908] = 0;
mem[909] = 0;
mem[910] = 1;
mem[911] = 1;
mem[912] = 1;
mem[913] = 1;
mem[914] = 0;
mem[915] = 0;
mem[916] = 0;
mem[917] = 0;
mem[918] = 0;
mem[919] = 0;
mem[920] = 0;
mem[921] = 0;
mem[922] = 0;
mem[923] = 0;
mem[924] = 0;
mem[925] = 0;
mem[926] = 1;
mem[927] = 1;
mem[928] = 1;
mem[929] = 1;
mem[930] = 1;
mem[931] = 0;
mem[932] = 0;
mem[933] = 0;
mem[934] = 0;
mem[935] = 0;
mem[936] = 0;
mem[937] = 0;
mem[938] = 0;
mem[939] = 1;
mem[940] = 1;
mem[941] = 1;
mem[942] = 0;
mem[943] = 0;
mem[944] = 0;
mem[945] = 0;
mem[946] = 0;
mem[947] = 0;
mem[948] = 0;
mem[949] = 0;
mem[950] = 0;
mem[951] = 0;
mem[952] = 0;
mem[953] = 0;
mem[954] = 0;
mem[955] = 0;
mem[956] = 0;
mem[957] = 0;
mem[958] = 0;
mem[959] = 0;
mem[960] = 0;
mem[961] = 1;
mem[962] = 1;
mem[963] = 0;
mem[964] = 0;
mem[965] = 0;
mem[966] = 0;
mem[967] = 0;
mem[968] = 0;
mem[969] = 0;
mem[970] = 0;
mem[971] = 0;
mem[972] = 1;
mem[973] = 1;
mem[974] = 1;
mem[975] = 1;
mem[976] = 1;
mem[977] = 0;
mem[978] = 0;
mem[979] = 0;
mem[980] = 1;
mem[981] = 1;
mem[982] = 0;
mem[983] = 0;
mem[984] = 0;
mem[985] = 0;
mem[986] = 0;
mem[987] = 0;
mem[988] = 0;
mem[989] = 0;
mem[990] = 0;
mem[991] = 0;
mem[992] = 0;
mem[993] = 0;
mem[994] = 1;
mem[995] = 1;
mem[996] = 1;
mem[997] = 1;
mem[998] = 1;
mem[999] = 1;
mem[1000] = 1;
mem[1001] = 1;
mem[1002] = 1;
mem[1003] = 1;
mem[1004] = 0;
mem[1005] = 0;
mem[1006] = 0;
mem[1007] = 0;
mem[1008] = 0;
mem[1009] = 0;
mem[1010] = 0;
mem[1011] = 0;
mem[1012] = 0;
mem[1013] = 0;
mem[1014] = 0;
mem[1015] = 0;
mem[1016] = 0;
mem[1017] = 1;
mem[1018] = 1;
mem[1019] = 1;
mem[1020] = 1;
mem[1021] = 0;
mem[1022] = 0;
mem[1023] = 0;
mem[1024] = 0;
mem[1025] = 0;
mem[1026] = 0;
mem[1027] = 0;
mem[1028] = 0;
mem[1029] = 1;
mem[1030] = 1;
mem[1031] = 0;
mem[1032] = 0;
mem[1033] = 0;
mem[1034] = 0;
mem[1035] = 0;
mem[1036] = 0;
mem[1037] = 0;
mem[1038] = 0;
mem[1039] = 0;
mem[1040] = 0;
mem[1041] = 0;
mem[1042] = 0;
mem[1043] = 0;
mem[1044] = 0;
mem[1045] = 0;
mem[1046] = 0;
mem[1047] = 0;
mem[1048] = 0;
mem[1049] = 0;
mem[1050] = 0;
mem[1051] = 0;
mem[1052] = 0;
mem[1053] = 0;
mem[1054] = 0;
mem[1055] = 0;
mem[1056] = 0;
mem[1057] = 0;
mem[1058] = 0;
mem[1059] = 0;
mem[1060] = 0;
mem[1061] = 0;
mem[1062] = 0;
mem[1063] = 1;
mem[1064] = 1;
mem[1065] = 0;
mem[1066] = 0;
mem[1067] = 0;
mem[1068] = 0;
mem[1069] = 0;
mem[1070] = 1;
mem[1071] = 1;
mem[1072] = 0;
mem[1073] = 0;
mem[1074] = 0;
mem[1075] = 0;
mem[1076] = 0;
mem[1077] = 0;
mem[1078] = 0;
mem[1079] = 0;
mem[1080] = 0;
mem[1081] = 1;
mem[1082] = 1;
mem[1083] = 1;
mem[1084] = 1;
mem[1085] = 1;
mem[1086] = 1;
mem[1087] = 1;
mem[1088] = 1;
mem[1089] = 1;
mem[1090] = 1;
mem[1091] = 0;
mem[1092] = 0;
mem[1093] = 0;
mem[1094] = 0;
mem[1095] = 0;
mem[1096] = 0;
mem[1097] = 0;
mem[1098] = 0;
mem[1099] = 0;
mem[1100] = 0;
mem[1101] = 0;
mem[1102] = 0;
mem[1103] = 0;
mem[1104] = 0;
mem[1105] = 0;
mem[1106] = 0;
mem[1107] = 0;
mem[1108] = 1;
mem[1109] = 1;
mem[1110] = 1;
mem[1111] = 0;
mem[1112] = 0;
mem[1113] = 0;
mem[1114] = 0;
mem[1115] = 0;
mem[1116] = 0;
mem[1117] = 0;
mem[1118] = 0;
mem[1119] = 0;
mem[1120] = 0;
mem[1121] = 0;
mem[1122] = 0;
mem[1123] = 0;
mem[1124] = 0;
mem[1125] = 0;
mem[1126] = 0;
mem[1127] = 0;
mem[1128] = 0;
mem[1129] = 0;
mem[1130] = 0;
mem[1131] = 0;
mem[1132] = 0;
mem[1133] = 0;
mem[1134] = 0;
mem[1135] = 0;
mem[1136] = 0;
mem[1137] = 0;
mem[1138] = 0;
mem[1139] = 0;
mem[1140] = 0;
mem[1141] = 0;
mem[1142] = 0;
mem[1143] = 0;
mem[1144] = 0;
mem[1145] = 0;
mem[1146] = 0;
mem[1147] = 0;
mem[1148] = 0;
mem[1149] = 0;
mem[1150] = 0;
mem[1151] = 0;
mem[1152] = 0;
mem[1153] = 0;
mem[1154] = 0;
mem[1155] = 0;
mem[1156] = 0;
mem[1157] = 0;
mem[1158] = 0;
mem[1159] = 0;
mem[1160] = 1;
mem[1161] = 1;
mem[1162] = 0;
mem[1163] = 0;
mem[1164] = 0;
mem[1165] = 0;
mem[1166] = 0;
mem[1167] = 0;
mem[1168] = 0;
mem[1169] = 0;
mem[1170] = 0;
mem[1171] = 1;
mem[1172] = 1;
mem[1173] = 1;
mem[1174] = 1;
mem[1175] = 1;
mem[1176] = 0;
mem[1177] = 0;
mem[1178] = 0;
mem[1179] = 0;
mem[1180] = 0;
mem[1181] = 0;
mem[1182] = 0;
mem[1183] = 0;
mem[1184] = 0;
mem[1185] = 0;
mem[1186] = 0;
mem[1187] = 0;
mem[1188] = 0;
mem[1189] = 0;
mem[1190] = 0;
mem[1191] = 0;
mem[1192] = 0;
mem[1193] = 0;
mem[1194] = 0;
mem[1195] = 0;
mem[1196] = 0;
mem[1197] = 0;
mem[1198] = 0;
mem[1199] = 0;
mem[1200] = 0;
mem[1201] = 0;
mem[1202] = 0;
mem[1203] = 0;
mem[1204] = 0;
mem[1205] = 0;
mem[1206] = 0;
mem[1207] = 0;
mem[1208] = 0;
mem[1209] = 0;
mem[1210] = 0;
mem[1211] = 0;
mem[1212] = 0;
mem[1213] = 0;
mem[1214] = 0;
mem[1215] = 0;
mem[1216] = 0;
mem[1217] = 0;
mem[1218] = 0;
mem[1219] = 0;
mem[1220] = 0;
mem[1221] = 0;
mem[1222] = 0;
mem[1223] = 0;
mem[1224] = 0;
mem[1225] = 0;
mem[1226] = 0;
mem[1227] = 0;
mem[1228] = 0;
mem[1229] = 0;
mem[1230] = 0;
mem[1231] = 0;
mem[1232] = 0;
mem[1233] = 0;
mem[1234] = 0;
mem[1235] = 0;
mem[1236] = 0;
mem[1237] = 0;
mem[1238] = 0;
mem[1239] = 0;
mem[1240] = 0;
mem[1241] = 0;
mem[1242] = 0;
mem[1243] = 0;
mem[1244] = 0;
mem[1245] = 0;
mem[1246] = 0;
mem[1247] = 0;
mem[1248] = 0;
mem[1249] = 1;
mem[1250] = 1;
mem[1251] = 1;
mem[1252] = 0;
mem[1253] = 0;
mem[1254] = 0;
mem[1255] = 0;
mem[1256] = 1;
mem[1257] = 1;
mem[1258] = 1;
mem[1259] = 1;
mem[1260] = 0;
mem[1261] = 0;
mem[1262] = 0;
mem[1263] = 1;
mem[1264] = 1;
mem[1265] = 1;
mem[1266] = 1;
mem[1267] = 1;
mem[1268] = 0;
mem[1269] = 0;
mem[1270] = 0;
mem[1271] = 0;
mem[1272] = 0;
mem[1273] = 0;
mem[1274] = 0;
mem[1275] = 0;
mem[1276] = 0;
mem[1277] = 0;
mem[1278] = 0;
mem[1279] = 0;
mem[1280] = 0;
mem[1281] = 0;
mem[1282] = 0;
mem[1283] = 0;
mem[1284] = 0;
mem[1285] = 0;
mem[1286] = 0;
mem[1287] = 0;
mem[1288] = 0;
mem[1289] = 0;
mem[1290] = 0;
mem[1291] = 0;
mem[1292] = 0;
mem[1293] = 0;
mem[1294] = 0;
mem[1295] = 0;
mem[1296] = 0;
mem[1297] = 0;
mem[1298] = 0;
mem[1299] = 0;
mem[1300] = 0;
mem[1301] = 0;
mem[1302] = 0;
mem[1303] = 0;
mem[1304] = 0;
mem[1305] = 0;
mem[1306] = 0;
mem[1307] = 0;
mem[1308] = 0;
mem[1309] = 0;
mem[1310] = 0;
mem[1311] = 0;
mem[1312] = 0;
mem[1313] = 0;
mem[1314] = 0;
mem[1315] = 0;
mem[1316] = 0;
mem[1317] = 0;
mem[1318] = 0;
mem[1319] = 0;
mem[1320] = 0;
mem[1321] = 0;
mem[1322] = 0;
mem[1323] = 0;
mem[1324] = 0;
mem[1325] = 0;
mem[1326] = 0;
mem[1327] = 0;
mem[1328] = 0;
mem[1329] = 0;
mem[1330] = 0;
mem[1331] = 0;
mem[1332] = 0;
mem[1333] = 0;
mem[1334] = 0;
mem[1335] = 0;
mem[1336] = 0;
mem[1337] = 0;
mem[1338] = 1;
mem[1339] = 1;
mem[1340] = 1;
mem[1341] = 1;
mem[1342] = 0;
mem[1343] = 0;
mem[1344] = 1;
mem[1345] = 1;
mem[1346] = 1;
mem[1347] = 1;
mem[1348] = 1;
mem[1349] = 1;
mem[1350] = 0;
mem[1351] = 0;
mem[1352] = 0;
mem[1353] = 0;
mem[1354] = 0;
mem[1355] = 1;
mem[1356] = 1;
mem[1357] = 1;
mem[1358] = 1;
mem[1359] = 1;
mem[1360] = 1;
mem[1361] = 0;
mem[1362] = 0;
mem[1363] = 0;
mem[1364] = 0;
mem[1365] = 0;
mem[1366] = 0;
mem[1367] = 0;
mem[1368] = 0;
mem[1369] = 0;
mem[1370] = 0;
mem[1371] = 0;
mem[1372] = 0;
mem[1373] = 0;
mem[1374] = 0;
mem[1375] = 0;
mem[1376] = 0;
mem[1377] = 0;
mem[1378] = 0;
mem[1379] = 0;
mem[1380] = 0;
mem[1381] = 0;
mem[1382] = 0;
mem[1383] = 0;
mem[1384] = 0;
mem[1385] = 0;
mem[1386] = 0;
mem[1387] = 0;
mem[1388] = 0;
mem[1389] = 0;
mem[1390] = 0;
mem[1391] = 0;
mem[1392] = 0;
mem[1393] = 0;
mem[1394] = 0;
mem[1395] = 0;
mem[1396] = 0;
mem[1397] = 0;
mem[1398] = 0;
mem[1399] = 0;
mem[1400] = 0;
mem[1401] = 0;
mem[1402] = 0;
mem[1403] = 0;
mem[1404] = 0;
mem[1405] = 0;
mem[1406] = 0;
mem[1407] = 0;
mem[1408] = 0;
mem[1409] = 0;
mem[1410] = 0;
mem[1411] = 0;
mem[1412] = 0;
mem[1413] = 0;
mem[1414] = 0;
mem[1415] = 0;
mem[1416] = 0;
mem[1417] = 0;
mem[1418] = 0;
mem[1419] = 0;
mem[1420] = 0;
mem[1421] = 0;
mem[1422] = 0;
mem[1423] = 0;
mem[1424] = 0;
mem[1425] = 0;
mem[1426] = 0;
mem[1427] = 0;
mem[1428] = 1;
mem[1429] = 1;
mem[1430] = 1;
mem[1431] = 1;
mem[1432] = 1;
mem[1433] = 1;
mem[1434] = 1;
mem[1435] = 1;
mem[1436] = 1;
mem[1437] = 1;
mem[1438] = 1;
mem[1439] = 1;
mem[1440] = 0;
mem[1441] = 0;
mem[1442] = 0;
mem[1443] = 0;
mem[1444] = 0;
mem[1445] = 0;
mem[1446] = 0;
mem[1447] = 1;
mem[1448] = 1;
mem[1449] = 1;
mem[1450] = 1;
mem[1451] = 1;
mem[1452] = 0;
mem[1453] = 0;
mem[1454] = 0;
mem[1455] = 0;
mem[1456] = 0;
mem[1457] = 0;
mem[1458] = 0;
mem[1459] = 0;
mem[1460] = 0;
mem[1461] = 0;
mem[1462] = 0;
mem[1463] = 0;
mem[1464] = 0;
mem[1465] = 0;
mem[1466] = 0;
mem[1467] = 0;
mem[1468] = 0;
mem[1469] = 0;
mem[1470] = 0;
mem[1471] = 0;
mem[1472] = 0;
mem[1473] = 0;
mem[1474] = 0;
mem[1475] = 0;
mem[1476] = 0;
mem[1477] = 0;
mem[1478] = 0;
mem[1479] = 0;
mem[1480] = 0;
mem[1481] = 0;
mem[1482] = 0;
mem[1483] = 0;
mem[1484] = 0;
mem[1485] = 0;
mem[1486] = 0;
mem[1487] = 0;
mem[1488] = 0;
mem[1489] = 0;
mem[1490] = 0;
mem[1491] = 0;
mem[1492] = 0;
mem[1493] = 0;
mem[1494] = 0;
mem[1495] = 0;
mem[1496] = 0;
mem[1497] = 0;
mem[1498] = 0;
mem[1499] = 0;
mem[1500] = 0;
mem[1501] = 0;
mem[1502] = 0;
mem[1503] = 0;
mem[1504] = 0;
mem[1505] = 0;
mem[1506] = 0;
mem[1507] = 0;
mem[1508] = 0;
mem[1509] = 0;
mem[1510] = 0;
mem[1511] = 0;
mem[1512] = 0;
mem[1513] = 0;
mem[1514] = 0;
mem[1515] = 0;
mem[1516] = 0;
mem[1517] = 0;
mem[1518] = 0;
mem[1519] = 1;
mem[1520] = 1;
mem[1521] = 1;
mem[1522] = 1;
mem[1523] = 1;
mem[1524] = 1;
mem[1525] = 1;
mem[1526] = 1;
mem[1527] = 1;
mem[1528] = 1;
mem[1529] = 1;
mem[1530] = 0;
mem[1531] = 0;
mem[1532] = 0;
mem[1533] = 0;
mem[1534] = 0;
mem[1535] = 0;
mem[1536] = 0;
mem[1537] = 0;
mem[1538] = 1;
mem[1539] = 1;
mem[1540] = 1;
mem[1541] = 1;
mem[1542] = 1;
mem[1543] = 0;
mem[1544] = 0;
mem[1545] = 0;
mem[1546] = 0;
mem[1547] = 0;
mem[1548] = 0;
mem[1549] = 0;
mem[1550] = 0;
mem[1551] = 0;
mem[1552] = 0;
mem[1553] = 0;
mem[1554] = 0;
mem[1555] = 0;
mem[1556] = 0;
mem[1557] = 0;
mem[1558] = 0;
mem[1559] = 0;
mem[1560] = 0;
mem[1561] = 0;
mem[1562] = 0;
mem[1563] = 0;
mem[1564] = 0;
mem[1565] = 0;
mem[1566] = 0;
mem[1567] = 0;
mem[1568] = 0;
mem[1569] = 0;
mem[1570] = 0;
mem[1571] = 0;
mem[1572] = 0;
mem[1573] = 0;
mem[1574] = 0;
mem[1575] = 0;
mem[1576] = 0;
mem[1577] = 0;
mem[1578] = 0;
mem[1579] = 0;
mem[1580] = 0;
mem[1581] = 0;
mem[1582] = 0;
mem[1583] = 0;
mem[1584] = 0;
mem[1585] = 0;
mem[1586] = 0;
mem[1587] = 0;
mem[1588] = 0;
mem[1589] = 0;
mem[1590] = 0;
mem[1591] = 0;
mem[1592] = 0;
mem[1593] = 0;
mem[1594] = 0;
mem[1595] = 0;
mem[1596] = 0;
mem[1597] = 0;
mem[1598] = 0;
mem[1599] = 0;
mem[1600] = 0;
mem[1601] = 0;
mem[1602] = 0;
mem[1603] = 0;
mem[1604] = 0;
mem[1605] = 0;
mem[1606] = 0;
mem[1607] = 0;
mem[1608] = 0;
mem[1609] = 0;
mem[1610] = 0;
mem[1611] = 0;
mem[1612] = 0;
mem[1613] = 0;
mem[1614] = 0;
mem[1615] = 1;
mem[1616] = 1;
mem[1617] = 1;
mem[1618] = 1;
mem[1619] = 0;
mem[1620] = 0;
mem[1621] = 0;
mem[1622] = 0;
mem[1623] = 0;
mem[1624] = 0;
mem[1625] = 0;
mem[1626] = 1;
mem[1627] = 1;
mem[1628] = 1;
mem[1629] = 1;
mem[1630] = 1;
mem[1631] = 1;
mem[1632] = 1;
mem[1633] = 0;
mem[1634] = 0;
mem[1635] = 0;
mem[1636] = 0;
mem[1637] = 0;
mem[1638] = 0;
mem[1639] = 0;
mem[1640] = 0;
mem[1641] = 0;
mem[1642] = 0;
mem[1643] = 0;
mem[1644] = 0;
mem[1645] = 0;
mem[1646] = 0;
mem[1647] = 0;
mem[1648] = 0;
mem[1649] = 0;
mem[1650] = 0;
mem[1651] = 0;
mem[1652] = 0;
mem[1653] = 0;
mem[1654] = 0;
mem[1655] = 0;
mem[1656] = 0;
mem[1657] = 0;
mem[1658] = 0;
mem[1659] = 0;
mem[1660] = 0;
mem[1661] = 0;
mem[1662] = 0;
mem[1663] = 0;
mem[1664] = 0;
mem[1665] = 0;
mem[1666] = 0;
mem[1667] = 0;
mem[1668] = 0;
mem[1669] = 0;
mem[1670] = 0;
mem[1671] = 0;
mem[1672] = 0;
mem[1673] = 0;
mem[1674] = 0;
mem[1675] = 0;
mem[1676] = 0;
mem[1677] = 0;
mem[1678] = 0;
mem[1679] = 0;
mem[1680] = 0;
mem[1681] = 0;
mem[1682] = 0;
mem[1683] = 0;
mem[1684] = 0;
mem[1685] = 0;
mem[1686] = 0;
mem[1687] = 0;
mem[1688] = 0;
mem[1689] = 0;
mem[1690] = 0;
mem[1691] = 0;
mem[1692] = 0;
mem[1693] = 0;
mem[1694] = 0;
mem[1695] = 0;
mem[1696] = 0;
mem[1697] = 0;
mem[1698] = 0;
mem[1699] = 0;
mem[1700] = 0;
mem[1701] = 0;
mem[1702] = 0;
mem[1703] = 0;
mem[1704] = 1;
mem[1705] = 1;
mem[1706] = 1;
mem[1707] = 0;
mem[1708] = 0;
mem[1709] = 0;
mem[1710] = 0;
mem[1711] = 1;
mem[1712] = 1;
mem[1713] = 1;
mem[1714] = 1;
mem[1715] = 1;
mem[1716] = 1;
mem[1717] = 1;
mem[1718] = 1;
mem[1719] = 1;
mem[1720] = 1;
mem[1721] = 0;
mem[1722] = 0;
mem[1723] = 0;
mem[1724] = 0;
mem[1725] = 0;
mem[1726] = 0;
mem[1727] = 0;
mem[1728] = 0;
mem[1729] = 0;
mem[1730] = 0;
mem[1731] = 0;
mem[1732] = 0;
mem[1733] = 0;
mem[1734] = 0;
mem[1735] = 0;
mem[1736] = 0;
mem[1737] = 0;
mem[1738] = 0;
mem[1739] = 0;
mem[1740] = 0;
mem[1741] = 0;
mem[1742] = 0;
mem[1743] = 0;
mem[1744] = 0;
mem[1745] = 0;
mem[1746] = 0;
mem[1747] = 0;
mem[1748] = 0;
mem[1749] = 0;
mem[1750] = 0;
mem[1751] = 0;
mem[1752] = 0;
mem[1753] = 0;
mem[1754] = 0;
mem[1755] = 0;
mem[1756] = 0;
mem[1757] = 0;
mem[1758] = 0;
mem[1759] = 0;
mem[1760] = 0;
mem[1761] = 0;
mem[1762] = 0;
mem[1763] = 0;
mem[1764] = 0;
mem[1765] = 0;
mem[1766] = 0;
mem[1767] = 0;
mem[1768] = 0;
mem[1769] = 0;
mem[1770] = 0;
mem[1771] = 0;
mem[1772] = 0;
mem[1773] = 0;
mem[1774] = 0;
mem[1775] = 0;
mem[1776] = 0;
mem[1777] = 0;
mem[1778] = 0;
mem[1779] = 0;
mem[1780] = 0;
mem[1781] = 0;
mem[1782] = 0;
mem[1783] = 0;
mem[1784] = 0;
mem[1785] = 0;
mem[1786] = 0;
mem[1787] = 0;
mem[1788] = 0;
mem[1789] = 0;
mem[1790] = 0;
mem[1791] = 1;
mem[1792] = 1;
mem[1793] = 1;
mem[1794] = 1;
mem[1795] = 1;
mem[1796] = 0;
mem[1797] = 0;
mem[1798] = 0;
mem[1799] = 0;
mem[1800] = 1;
mem[1801] = 1;
mem[1802] = 1;
mem[1803] = 1;
mem[1804] = 1;
mem[1805] = 1;
mem[1806] = 1;
mem[1807] = 1;
mem[1808] = 1;
mem[1809] = 0;
mem[1810] = 0;
mem[1811] = 0;
mem[1812] = 0;
mem[1813] = 0;
mem[1814] = 0;
mem[1815] = 0;
mem[1816] = 0;
mem[1817] = 0;
mem[1818] = 0;
mem[1819] = 0;
mem[1820] = 0;
mem[1821] = 0;
mem[1822] = 0;
mem[1823] = 0;
mem[1824] = 0;
mem[1825] = 0;
mem[1826] = 0;
mem[1827] = 0;
mem[1828] = 0;
mem[1829] = 0;
mem[1830] = 0;
mem[1831] = 0;
mem[1832] = 0;
mem[1833] = 0;
mem[1834] = 0;
mem[1835] = 0;
mem[1836] = 0;
mem[1837] = 0;
mem[1838] = 0;
mem[1839] = 0;
mem[1840] = 0;
mem[1841] = 0;
mem[1842] = 0;
mem[1843] = 0;
mem[1844] = 0;
mem[1845] = 0;
mem[1846] = 0;
mem[1847] = 0;
mem[1848] = 0;
mem[1849] = 0;
mem[1850] = 0;
mem[1851] = 0;
mem[1852] = 0;
mem[1853] = 0;
mem[1854] = 0;
mem[1855] = 0;
mem[1856] = 0;
mem[1857] = 0;
mem[1858] = 0;
mem[1859] = 0;
mem[1860] = 0;
mem[1861] = 0;
mem[1862] = 0;
mem[1863] = 0;
mem[1864] = 0;
mem[1865] = 0;
mem[1866] = 0;
mem[1867] = 0;
mem[1868] = 0;
mem[1869] = 0;
mem[1870] = 0;
mem[1871] = 0;
mem[1872] = 0;
mem[1873] = 0;
mem[1874] = 0;
mem[1875] = 0;
mem[1876] = 0;
mem[1877] = 0;
mem[1878] = 0;
mem[1879] = 0;
mem[1880] = 1;
mem[1881] = 1;
mem[1882] = 1;
mem[1883] = 1;
mem[1884] = 1;
mem[1885] = 0;
mem[1886] = 0;
mem[1887] = 0;
mem[1888] = 0;
mem[1889] = 0;
mem[1890] = 1;
mem[1891] = 1;
mem[1892] = 1;
mem[1893] = 1;
mem[1894] = 1;
mem[1895] = 1;
mem[1896] = 0;
mem[1897] = 0;
mem[1898] = 0;
mem[1899] = 0;
mem[1900] = 0;
mem[1901] = 0;
mem[1902] = 0;
mem[1903] = 0;
mem[1904] = 0;
mem[1905] = 0;
mem[1906] = 0;
mem[1907] = 0;
mem[1908] = 0;
mem[1909] = 0;
mem[1910] = 0;
mem[1911] = 0;
mem[1912] = 0;
mem[1913] = 0;
mem[1914] = 0;
mem[1915] = 0;
mem[1916] = 0;
mem[1917] = 0;
mem[1918] = 0;
mem[1919] = 0;
mem[1920] = 0;
mem[1921] = 0;
mem[1922] = 0;
mem[1923] = 0;
mem[1924] = 0;
mem[1925] = 0;
mem[1926] = 0;
mem[1927] = 0;
mem[1928] = 0;
mem[1929] = 0;
mem[1930] = 0;
mem[1931] = 0;
mem[1932] = 0;
mem[1933] = 0;
mem[1934] = 0;
mem[1935] = 0;
mem[1936] = 0;
mem[1937] = 0;
mem[1938] = 0;
mem[1939] = 0;
mem[1940] = 0;
mem[1941] = 0;
mem[1942] = 0;
mem[1943] = 0;
mem[1944] = 0;
mem[1945] = 0;
mem[1946] = 0;
mem[1947] = 0;
mem[1948] = 0;
mem[1949] = 0;
mem[1950] = 0;
mem[1951] = 0;
mem[1952] = 0;
mem[1953] = 0;
mem[1954] = 0;
mem[1955] = 0;
mem[1956] = 0;
mem[1957] = 0;
mem[1958] = 0;
mem[1959] = 0;
mem[1960] = 0;
mem[1961] = 0;
mem[1962] = 0;
mem[1963] = 0;
mem[1964] = 0;
mem[1965] = 0;
mem[1966] = 0;
mem[1967] = 0;
mem[1968] = 0;
mem[1969] = 0;
mem[1970] = 1;
mem[1971] = 1;
mem[1972] = 1;
mem[1973] = 0;
mem[1974] = 0;
mem[1975] = 0;
mem[1976] = 0;
mem[1977] = 0;
mem[1978] = 0;
mem[1979] = 0;
mem[1980] = 1;
mem[1981] = 1;
mem[1982] = 1;
mem[1983] = 0;
mem[1984] = 0;
mem[1985] = 0;
mem[1986] = 0;
mem[1987] = 0;
mem[1988] = 0;
mem[1989] = 0;
mem[1990] = 0;
mem[1991] = 0;
mem[1992] = 0;
mem[1993] = 0;
mem[1994] = 0;
mem[1995] = 0;
mem[1996] = 0;
mem[1997] = 0;
mem[1998] = 0;
mem[1999] = 1;
mem[2000] = 1;
mem[2001] = 0;
mem[2002] = 0;
mem[2003] = 0;
mem[2004] = 0;
mem[2005] = 1;
mem[2006] = 1;
mem[2007] = 0;
mem[2008] = 0;
mem[2009] = 1;
mem[2010] = 1;
mem[2011] = 1;
mem[2012] = 1;
mem[2013] = 0;
mem[2014] = 0;
mem[2015] = 1;
mem[2016] = 1;
mem[2017] = 0;
mem[2018] = 0;
mem[2019] = 0;
mem[2020] = 0;
mem[2021] = 1;
mem[2022] = 1;
mem[2023] = 0;
mem[2024] = 0;
mem[2025] = 1;
mem[2026] = 1;
mem[2027] = 0;
mem[2028] = 0;
mem[2029] = 0;
mem[2030] = 0;
mem[2031] = 1;
mem[2032] = 1;
mem[2033] = 0;
mem[2034] = 1;
mem[2035] = 1;
mem[2036] = 1;
mem[2037] = 1;
mem[2038] = 1;
mem[2039] = 1;
mem[2040] = 1;
mem[2041] = 0;
mem[2042] = 0;
mem[2043] = 1;
mem[2044] = 1;
mem[2045] = 1;
mem[2046] = 1;
mem[2047] = 1;
mem[2048] = 1;
mem[2049] = 0;
mem[2050] = 0;
mem[2051] = 0;
mem[2052] = 0;
mem[2053] = 0;
mem[2054] = 0;
mem[2055] = 0;
mem[2056] = 0;
mem[2057] = 0;
mem[2058] = 0;
mem[2059] = 0;
mem[2060] = 1;
mem[2061] = 1;
mem[2062] = 1;
mem[2063] = 0;
mem[2064] = 0;
mem[2065] = 0;
mem[2066] = 0;
mem[2067] = 0;
mem[2068] = 0;
mem[2069] = 0;
mem[2070] = 1;
mem[2071] = 1;
mem[2072] = 1;
mem[2073] = 1;
mem[2074] = 1;
mem[2075] = 1;
mem[2076] = 0;
mem[2077] = 0;
mem[2078] = 0;
mem[2079] = 0;
mem[2080] = 0;
mem[2081] = 0;
mem[2082] = 0;
mem[2083] = 0;
mem[2084] = 0;
mem[2085] = 0;
mem[2086] = 0;
mem[2087] = 0;
mem[2088] = 0;
mem[2089] = 1;
mem[2090] = 1;
mem[2091] = 0;
mem[2092] = 0;
mem[2093] = 0;
mem[2094] = 0;
mem[2095] = 1;
mem[2096] = 1;
mem[2097] = 0;
mem[2098] = 0;
mem[2099] = 1;
mem[2100] = 1;
mem[2101] = 1;
mem[2102] = 1;
mem[2103] = 0;
mem[2104] = 0;
mem[2105] = 1;
mem[2106] = 1;
mem[2107] = 0;
mem[2108] = 0;
mem[2109] = 0;
mem[2110] = 0;
mem[2111] = 1;
mem[2112] = 1;
mem[2113] = 0;
mem[2114] = 0;
mem[2115] = 1;
mem[2116] = 1;
mem[2117] = 0;
mem[2118] = 0;
mem[2119] = 0;
mem[2120] = 0;
mem[2121] = 1;
mem[2122] = 1;
mem[2123] = 0;
mem[2124] = 1;
mem[2125] = 1;
mem[2126] = 1;
mem[2127] = 1;
mem[2128] = 1;
mem[2129] = 1;
mem[2130] = 1;
mem[2131] = 0;
mem[2132] = 0;
mem[2133] = 1;
mem[2134] = 1;
mem[2135] = 1;
mem[2136] = 1;
mem[2137] = 1;
mem[2138] = 1;
mem[2139] = 1;
mem[2140] = 0;
mem[2141] = 0;
mem[2142] = 0;
mem[2143] = 0;
mem[2144] = 0;
mem[2145] = 0;
mem[2146] = 0;
mem[2147] = 0;
mem[2148] = 0;
mem[2149] = 0;
mem[2150] = 1;
mem[2151] = 1;
mem[2152] = 1;
mem[2153] = 1;
mem[2154] = 1;
mem[2155] = 0;
mem[2156] = 0;
mem[2157] = 0;
mem[2158] = 0;
mem[2159] = 0;
mem[2160] = 0;
mem[2161] = 0;
mem[2162] = 1;
mem[2163] = 1;
mem[2164] = 1;
mem[2165] = 1;
mem[2166] = 1;
mem[2167] = 1;
mem[2168] = 1;
mem[2169] = 0;
mem[2170] = 0;
mem[2171] = 0;
mem[2172] = 0;
mem[2173] = 0;
mem[2174] = 0;
mem[2175] = 0;
mem[2176] = 0;
mem[2177] = 0;
mem[2178] = 0;
mem[2179] = 1;
mem[2180] = 1;
mem[2181] = 0;
mem[2182] = 0;
mem[2183] = 0;
mem[2184] = 0;
mem[2185] = 1;
mem[2186] = 1;
mem[2187] = 0;
mem[2188] = 0;
mem[2189] = 0;
mem[2190] = 1;
mem[2191] = 1;
mem[2192] = 0;
mem[2193] = 0;
mem[2194] = 0;
mem[2195] = 1;
mem[2196] = 1;
mem[2197] = 1;
mem[2198] = 0;
mem[2199] = 0;
mem[2200] = 0;
mem[2201] = 1;
mem[2202] = 1;
mem[2203] = 0;
mem[2204] = 0;
mem[2205] = 1;
mem[2206] = 1;
mem[2207] = 1;
mem[2208] = 0;
mem[2209] = 0;
mem[2210] = 0;
mem[2211] = 1;
mem[2212] = 1;
mem[2213] = 0;
mem[2214] = 1;
mem[2215] = 1;
mem[2216] = 0;
mem[2217] = 0;
mem[2218] = 0;
mem[2219] = 0;
mem[2220] = 0;
mem[2221] = 0;
mem[2222] = 0;
mem[2223] = 1;
mem[2224] = 1;
mem[2225] = 0;
mem[2226] = 0;
mem[2227] = 1;
mem[2228] = 1;
mem[2229] = 1;
mem[2230] = 0;
mem[2231] = 0;
mem[2232] = 0;
mem[2233] = 0;
mem[2234] = 0;
mem[2235] = 0;
mem[2236] = 0;
mem[2237] = 0;
mem[2238] = 0;
mem[2239] = 0;
mem[2240] = 0;
mem[2241] = 0;
mem[2242] = 1;
mem[2243] = 1;
mem[2244] = 1;
mem[2245] = 1;
mem[2246] = 1;
mem[2247] = 0;
mem[2248] = 0;
mem[2249] = 0;
mem[2250] = 0;
mem[2251] = 0;
mem[2252] = 0;
mem[2253] = 0;
mem[2254] = 0;
mem[2255] = 0;
mem[2256] = 1;
mem[2257] = 1;
mem[2258] = 1;
mem[2259] = 1;
mem[2260] = 1;
mem[2261] = 0;
mem[2262] = 0;
mem[2263] = 0;
mem[2264] = 0;
mem[2265] = 0;
mem[2266] = 0;
mem[2267] = 0;
mem[2268] = 0;
mem[2269] = 1;
mem[2270] = 1;
mem[2271] = 0;
mem[2272] = 0;
mem[2273] = 0;
mem[2274] = 0;
mem[2275] = 1;
mem[2276] = 1;
mem[2277] = 0;
mem[2278] = 0;
mem[2279] = 0;
mem[2280] = 1;
mem[2281] = 1;
mem[2282] = 0;
mem[2283] = 0;
mem[2284] = 0;
mem[2285] = 1;
mem[2286] = 1;
mem[2287] = 1;
mem[2288] = 1;
mem[2289] = 0;
mem[2290] = 0;
mem[2291] = 1;
mem[2292] = 1;
mem[2293] = 0;
mem[2294] = 0;
mem[2295] = 1;
mem[2296] = 1;
mem[2297] = 1;
mem[2298] = 1;
mem[2299] = 0;
mem[2300] = 0;
mem[2301] = 1;
mem[2302] = 1;
mem[2303] = 0;
mem[2304] = 1;
mem[2305] = 1;
mem[2306] = 0;
mem[2307] = 0;
mem[2308] = 0;
mem[2309] = 0;
mem[2310] = 0;
mem[2311] = 0;
mem[2312] = 0;
mem[2313] = 1;
mem[2314] = 1;
mem[2315] = 0;
mem[2316] = 0;
mem[2317] = 1;
mem[2318] = 1;
mem[2319] = 1;
mem[2320] = 0;
mem[2321] = 0;
mem[2322] = 0;
mem[2323] = 0;
mem[2324] = 0;
mem[2325] = 0;
mem[2326] = 0;
mem[2327] = 0;
mem[2328] = 0;
mem[2329] = 0;
mem[2330] = 0;
mem[2331] = 0;
mem[2332] = 0;
mem[2333] = 0;
mem[2334] = 0;
mem[2335] = 1;
mem[2336] = 1;
mem[2337] = 1;
mem[2338] = 0;
mem[2339] = 0;
mem[2340] = 0;
mem[2341] = 0;
mem[2342] = 0;
mem[2343] = 0;
mem[2344] = 0;
mem[2345] = 0;
mem[2346] = 0;
mem[2347] = 0;
mem[2348] = 1;
mem[2349] = 1;
mem[2350] = 1;
mem[2351] = 1;
mem[2352] = 0;
mem[2353] = 0;
mem[2354] = 0;
mem[2355] = 0;
mem[2356] = 0;
mem[2357] = 0;
mem[2358] = 0;
mem[2359] = 1;
mem[2360] = 1;
mem[2361] = 0;
mem[2362] = 1;
mem[2363] = 1;
mem[2364] = 0;
mem[2365] = 1;
mem[2366] = 1;
mem[2367] = 0;
mem[2368] = 0;
mem[2369] = 0;
mem[2370] = 1;
mem[2371] = 1;
mem[2372] = 0;
mem[2373] = 0;
mem[2374] = 0;
mem[2375] = 1;
mem[2376] = 1;
mem[2377] = 1;
mem[2378] = 1;
mem[2379] = 1;
mem[2380] = 0;
mem[2381] = 1;
mem[2382] = 1;
mem[2383] = 0;
mem[2384] = 0;
mem[2385] = 1;
mem[2386] = 1;
mem[2387] = 1;
mem[2388] = 1;
mem[2389] = 1;
mem[2390] = 0;
mem[2391] = 1;
mem[2392] = 1;
mem[2393] = 0;
mem[2394] = 1;
mem[2395] = 1;
mem[2396] = 0;
mem[2397] = 0;
mem[2398] = 0;
mem[2399] = 0;
mem[2400] = 0;
mem[2401] = 0;
mem[2402] = 0;
mem[2403] = 1;
mem[2404] = 1;
mem[2405] = 0;
mem[2406] = 0;
mem[2407] = 1;
mem[2408] = 1;
mem[2409] = 1;
mem[2410] = 0;
mem[2411] = 0;
mem[2412] = 0;
mem[2413] = 0;
mem[2414] = 0;
mem[2415] = 0;
mem[2416] = 0;
mem[2417] = 0;
mem[2418] = 0;
mem[2419] = 0;
mem[2420] = 0;
mem[2421] = 0;
mem[2422] = 0;
mem[2423] = 0;
mem[2424] = 0;
mem[2425] = 0;
mem[2426] = 0;
mem[2427] = 1;
mem[2428] = 1;
mem[2429] = 1;
mem[2430] = 0;
mem[2431] = 0;
mem[2432] = 0;
mem[2433] = 0;
mem[2434] = 0;
mem[2435] = 1;
mem[2436] = 1;
mem[2437] = 1;
mem[2438] = 1;
mem[2439] = 1;
mem[2440] = 0;
mem[2441] = 0;
mem[2442] = 0;
mem[2443] = 0;
mem[2444] = 0;
mem[2445] = 0;
mem[2446] = 0;
mem[2447] = 0;
mem[2448] = 0;
mem[2449] = 1;
mem[2450] = 1;
mem[2451] = 0;
mem[2452] = 1;
mem[2453] = 1;
mem[2454] = 0;
mem[2455] = 1;
mem[2456] = 1;
mem[2457] = 0;
mem[2458] = 0;
mem[2459] = 0;
mem[2460] = 1;
mem[2461] = 1;
mem[2462] = 0;
mem[2463] = 0;
mem[2464] = 0;
mem[2465] = 1;
mem[2466] = 1;
mem[2467] = 0;
mem[2468] = 1;
mem[2469] = 1;
mem[2470] = 1;
mem[2471] = 1;
mem[2472] = 1;
mem[2473] = 0;
mem[2474] = 0;
mem[2475] = 1;
mem[2476] = 1;
mem[2477] = 0;
mem[2478] = 1;
mem[2479] = 1;
mem[2480] = 1;
mem[2481] = 1;
mem[2482] = 1;
mem[2483] = 0;
mem[2484] = 1;
mem[2485] = 1;
mem[2486] = 1;
mem[2487] = 1;
mem[2488] = 1;
mem[2489] = 1;
mem[2490] = 1;
mem[2491] = 0;
mem[2492] = 0;
mem[2493] = 1;
mem[2494] = 1;
mem[2495] = 1;
mem[2496] = 1;
mem[2497] = 1;
mem[2498] = 1;
mem[2499] = 0;
mem[2500] = 0;
mem[2501] = 0;
mem[2502] = 0;
mem[2503] = 0;
mem[2504] = 0;
mem[2505] = 0;
mem[2506] = 0;
mem[2507] = 0;
mem[2508] = 0;
mem[2509] = 0;
mem[2510] = 0;
mem[2511] = 0;
mem[2512] = 0;
mem[2513] = 0;
mem[2514] = 0;
mem[2515] = 0;
mem[2516] = 0;
mem[2517] = 1;
mem[2518] = 1;
mem[2519] = 1;
mem[2520] = 0;
mem[2521] = 0;
mem[2522] = 0;
mem[2523] = 1;
mem[2524] = 1;
mem[2525] = 1;
mem[2526] = 1;
mem[2527] = 1;
mem[2528] = 0;
mem[2529] = 0;
mem[2530] = 0;
mem[2531] = 0;
mem[2532] = 0;
mem[2533] = 0;
mem[2534] = 0;
mem[2535] = 0;
mem[2536] = 0;
mem[2537] = 0;
mem[2538] = 0;
mem[2539] = 1;
mem[2540] = 1;
mem[2541] = 0;
mem[2542] = 1;
mem[2543] = 1;
mem[2544] = 0;
mem[2545] = 1;
mem[2546] = 1;
mem[2547] = 0;
mem[2548] = 0;
mem[2549] = 0;
mem[2550] = 1;
mem[2551] = 1;
mem[2552] = 0;
mem[2553] = 0;
mem[2554] = 0;
mem[2555] = 1;
mem[2556] = 1;
mem[2557] = 0;
mem[2558] = 0;
mem[2559] = 1;
mem[2560] = 1;
mem[2561] = 1;
mem[2562] = 1;
mem[2563] = 0;
mem[2564] = 0;
mem[2565] = 1;
mem[2566] = 1;
mem[2567] = 0;
mem[2568] = 0;
mem[2569] = 1;
mem[2570] = 1;
mem[2571] = 1;
mem[2572] = 1;
mem[2573] = 0;
mem[2574] = 1;
mem[2575] = 1;
mem[2576] = 1;
mem[2577] = 1;
mem[2578] = 1;
mem[2579] = 1;
mem[2580] = 1;
mem[2581] = 0;
mem[2582] = 0;
mem[2583] = 1;
mem[2584] = 1;
mem[2585] = 1;
mem[2586] = 1;
mem[2587] = 1;
mem[2588] = 1;
mem[2589] = 0;
mem[2590] = 0;
mem[2591] = 0;
mem[2592] = 0;
mem[2593] = 0;
mem[2594] = 0;
mem[2595] = 0;
mem[2596] = 0;
mem[2597] = 0;
mem[2598] = 0;
mem[2599] = 0;
mem[2600] = 0;
mem[2601] = 0;
mem[2602] = 0;
mem[2603] = 0;
mem[2604] = 1;
mem[2605] = 1;
mem[2606] = 1;
mem[2607] = 1;
mem[2608] = 0;
mem[2609] = 0;
mem[2610] = 0;
mem[2611] = 1;
mem[2612] = 1;
mem[2613] = 1;
mem[2614] = 1;
mem[2615] = 1;
mem[2616] = 0;
mem[2617] = 0;
mem[2618] = 0;
mem[2619] = 0;
mem[2620] = 0;
mem[2621] = 0;
mem[2622] = 0;
mem[2623] = 0;
mem[2624] = 0;
mem[2625] = 0;
mem[2626] = 0;
mem[2627] = 0;
mem[2628] = 0;
mem[2629] = 1;
mem[2630] = 1;
mem[2631] = 1;
mem[2632] = 1;
mem[2633] = 1;
mem[2634] = 1;
mem[2635] = 1;
mem[2636] = 1;
mem[2637] = 0;
mem[2638] = 0;
mem[2639] = 0;
mem[2640] = 1;
mem[2641] = 1;
mem[2642] = 0;
mem[2643] = 0;
mem[2644] = 0;
mem[2645] = 1;
mem[2646] = 1;
mem[2647] = 0;
mem[2648] = 0;
mem[2649] = 0;
mem[2650] = 1;
mem[2651] = 1;
mem[2652] = 1;
mem[2653] = 0;
mem[2654] = 0;
mem[2655] = 1;
mem[2656] = 1;
mem[2657] = 0;
mem[2658] = 0;
mem[2659] = 0;
mem[2660] = 1;
mem[2661] = 1;
mem[2662] = 1;
mem[2663] = 0;
mem[2664] = 1;
mem[2665] = 1;
mem[2666] = 0;
mem[2667] = 0;
mem[2668] = 0;
mem[2669] = 0;
mem[2670] = 0;
mem[2671] = 0;
mem[2672] = 0;
mem[2673] = 1;
mem[2674] = 1;
mem[2675] = 0;
mem[2676] = 1;
mem[2677] = 1;
mem[2678] = 1;
mem[2679] = 1;
mem[2680] = 0;
mem[2681] = 0;
mem[2682] = 0;
mem[2683] = 0;
mem[2684] = 0;
mem[2685] = 0;
mem[2686] = 0;
mem[2687] = 0;
mem[2688] = 0;
mem[2689] = 0;
mem[2690] = 0;
mem[2691] = 1;
mem[2692] = 1;
mem[2693] = 1;
mem[2694] = 1;
mem[2695] = 1;
mem[2696] = 1;
mem[2697] = 0;
mem[2698] = 0;
mem[2699] = 0;
mem[2700] = 0;
mem[2701] = 1;
mem[2702] = 1;
mem[2703] = 1;
mem[2704] = 0;
mem[2705] = 0;
mem[2706] = 0;
mem[2707] = 0;
mem[2708] = 0;
mem[2709] = 0;
mem[2710] = 0;
mem[2711] = 0;
mem[2712] = 0;
mem[2713] = 0;
mem[2714] = 0;
mem[2715] = 0;
mem[2716] = 0;
mem[2717] = 0;
mem[2718] = 0;
mem[2719] = 0;
mem[2720] = 1;
mem[2721] = 1;
mem[2722] = 0;
mem[2723] = 0;
mem[2724] = 1;
mem[2725] = 1;
mem[2726] = 0;
mem[2727] = 0;
mem[2728] = 0;
mem[2729] = 0;
mem[2730] = 1;
mem[2731] = 1;
mem[2732] = 0;
mem[2733] = 0;
mem[2734] = 0;
mem[2735] = 1;
mem[2736] = 1;
mem[2737] = 0;
mem[2738] = 0;
mem[2739] = 0;
mem[2740] = 0;
mem[2741] = 1;
mem[2742] = 1;
mem[2743] = 0;
mem[2744] = 0;
mem[2745] = 1;
mem[2746] = 1;
mem[2747] = 0;
mem[2748] = 0;
mem[2749] = 0;
mem[2750] = 0;
mem[2751] = 1;
mem[2752] = 1;
mem[2753] = 0;
mem[2754] = 1;
mem[2755] = 1;
mem[2756] = 0;
mem[2757] = 0;
mem[2758] = 0;
mem[2759] = 0;
mem[2760] = 0;
mem[2761] = 0;
mem[2762] = 0;
mem[2763] = 1;
mem[2764] = 1;
mem[2765] = 0;
mem[2766] = 0;
mem[2767] = 1;
mem[2768] = 1;
mem[2769] = 1;
mem[2770] = 0;
mem[2771] = 0;
mem[2772] = 0;
mem[2773] = 0;
mem[2774] = 0;
mem[2775] = 0;
mem[2776] = 0;
mem[2777] = 0;
mem[2778] = 0;
mem[2779] = 0;
mem[2780] = 1;
mem[2781] = 1;
mem[2782] = 1;
mem[2783] = 1;
mem[2784] = 0;
mem[2785] = 0;
mem[2786] = 0;
mem[2787] = 0;
mem[2788] = 0;
mem[2789] = 0;
mem[2790] = 0;
mem[2791] = 1;
mem[2792] = 1;
mem[2793] = 1;
mem[2794] = 1;
mem[2795] = 1;
mem[2796] = 0;
mem[2797] = 0;
mem[2798] = 0;
mem[2799] = 0;
mem[2800] = 0;
mem[2801] = 0;
mem[2802] = 0;
mem[2803] = 0;
mem[2804] = 0;
mem[2805] = 0;
mem[2806] = 0;
mem[2807] = 0;
mem[2808] = 0;
mem[2809] = 0;
mem[2810] = 1;
mem[2811] = 1;
mem[2812] = 0;
mem[2813] = 0;
mem[2814] = 1;
mem[2815] = 1;
mem[2816] = 0;
mem[2817] = 0;
mem[2818] = 0;
mem[2819] = 1;
mem[2820] = 1;
mem[2821] = 1;
mem[2822] = 1;
mem[2823] = 0;
mem[2824] = 0;
mem[2825] = 1;
mem[2826] = 1;
mem[2827] = 0;
mem[2828] = 0;
mem[2829] = 0;
mem[2830] = 0;
mem[2831] = 1;
mem[2832] = 1;
mem[2833] = 0;
mem[2834] = 0;
mem[2835] = 1;
mem[2836] = 1;
mem[2837] = 0;
mem[2838] = 0;
mem[2839] = 0;
mem[2840] = 0;
mem[2841] = 1;
mem[2842] = 1;
mem[2843] = 0;
mem[2844] = 1;
mem[2845] = 1;
mem[2846] = 1;
mem[2847] = 1;
mem[2848] = 1;
mem[2849] = 1;
mem[2850] = 1;
mem[2851] = 0;
mem[2852] = 0;
mem[2853] = 1;
mem[2854] = 1;
mem[2855] = 0;
mem[2856] = 0;
mem[2857] = 0;
mem[2858] = 1;
mem[2859] = 1;
mem[2860] = 0;
mem[2861] = 0;
mem[2862] = 0;
mem[2863] = 0;
mem[2864] = 0;
mem[2865] = 0;
mem[2866] = 0;
mem[2867] = 0;
mem[2868] = 0;
mem[2869] = 1;
mem[2870] = 1;
mem[2871] = 1;
mem[2872] = 0;
mem[2873] = 0;
mem[2874] = 0;
mem[2875] = 0;
mem[2876] = 0;
mem[2877] = 0;
mem[2878] = 0;
mem[2879] = 0;
mem[2880] = 0;
mem[2881] = 0;
mem[2882] = 0;
mem[2883] = 1;
mem[2884] = 1;
mem[2885] = 1;
mem[2886] = 1;
mem[2887] = 1;
mem[2888] = 0;
mem[2889] = 0;
mem[2890] = 0;
mem[2891] = 0;
mem[2892] = 0;
mem[2893] = 0;
mem[2894] = 0;
mem[2895] = 0;
mem[2896] = 0;
mem[2897] = 0;
mem[2898] = 0;
mem[2899] = 0;
mem[2900] = 1;
mem[2901] = 1;
mem[2902] = 0;
mem[2903] = 0;
mem[2904] = 1;
mem[2905] = 1;
mem[2906] = 0;
mem[2907] = 0;
mem[2908] = 0;
mem[2909] = 1;
mem[2910] = 1;
mem[2911] = 1;
mem[2912] = 1;
mem[2913] = 0;
mem[2914] = 0;
mem[2915] = 1;
mem[2916] = 1;
mem[2917] = 0;
mem[2918] = 0;
mem[2919] = 0;
mem[2920] = 0;
mem[2921] = 1;
mem[2922] = 1;
mem[2923] = 0;
mem[2924] = 0;
mem[2925] = 1;
mem[2926] = 1;
mem[2927] = 0;
mem[2928] = 0;
mem[2929] = 0;
mem[2930] = 0;
mem[2931] = 1;
mem[2932] = 1;
mem[2933] = 0;
mem[2934] = 1;
mem[2935] = 1;
mem[2936] = 1;
mem[2937] = 1;
mem[2938] = 1;
mem[2939] = 1;
mem[2940] = 1;
mem[2941] = 0;
mem[2942] = 0;
mem[2943] = 1;
mem[2944] = 1;
mem[2945] = 0;
mem[2946] = 0;
mem[2947] = 0;
mem[2948] = 1;
mem[2949] = 1;
mem[2950] = 0;
mem[2951] = 0;
mem[2952] = 0;
mem[2953] = 0;
mem[2954] = 0;
mem[2955] = 0;
mem[2956] = 0;
mem[2957] = 0;
mem[2958] = 0;
mem[2959] = 1;
mem[2960] = 1;
mem[2961] = 1;
mem[2962] = 0;
mem[2963] = 0;
mem[2964] = 0;
mem[2965] = 0;
mem[2966] = 0;
mem[2967] = 0;
mem[2968] = 0;
mem[2969] = 0;
mem[2970] = 0;
mem[2971] = 0;
mem[2972] = 0;
mem[2973] = 0;
mem[2974] = 0;
mem[2975] = 1;
mem[2976] = 1;
mem[2977] = 1;
mem[2978] = 1;
mem[2979] = 1;
mem[2980] = 1;
mem[2981] = 0;
mem[2982] = 0;
mem[2983] = 0;
mem[2984] = 0;
mem[2985] = 0;
mem[2986] = 0;
mem[2987] = 0;
mem[2988] = 0;
mem[2989] = 0;
mem[2990] = 0;
mem[2991] = 0;
mem[2992] = 0;
mem[2993] = 0;
mem[2994] = 0;
mem[2995] = 0;
mem[2996] = 0;
mem[2997] = 0;
mem[2998] = 0;
mem[2999] = 0;
mem[3000] = 0;
mem[3001] = 0;
mem[3002] = 0;
mem[3003] = 0;
mem[3004] = 0;
mem[3005] = 0;
mem[3006] = 0;
mem[3007] = 0;
mem[3008] = 0;
mem[3009] = 0;
mem[3010] = 0;
mem[3011] = 0;
mem[3012] = 0;
mem[3013] = 0;
mem[3014] = 0;
mem[3015] = 0;
mem[3016] = 0;
mem[3017] = 0;
mem[3018] = 0;
mem[3019] = 0;
mem[3020] = 0;
mem[3021] = 0;
mem[3022] = 0;
mem[3023] = 0;
mem[3024] = 0;
mem[3025] = 0;
mem[3026] = 0;
mem[3027] = 0;
mem[3028] = 0;
mem[3029] = 0;
mem[3030] = 0;
mem[3031] = 0;
mem[3032] = 0;
mem[3033] = 0;
mem[3034] = 0;
mem[3035] = 0;
mem[3036] = 0;
mem[3037] = 0;
mem[3038] = 0;
mem[3039] = 0;
mem[3040] = 0;
mem[3041] = 0;
mem[3042] = 0;
mem[3043] = 0;
mem[3044] = 0;
mem[3045] = 0;
mem[3046] = 0;
mem[3047] = 0;
mem[3048] = 0;
mem[3049] = 1;
mem[3050] = 1;
mem[3051] = 1;
mem[3052] = 1;
mem[3053] = 0;
mem[3054] = 0;
mem[3055] = 0;
mem[3056] = 0;
mem[3057] = 0;
mem[3058] = 0;
mem[3059] = 0;
mem[3060] = 0;
mem[3061] = 0;
mem[3062] = 0;
mem[3063] = 0;
mem[3064] = 0;
mem[3065] = 0;
mem[3066] = 1;
mem[3067] = 1;
mem[3068] = 1;
mem[3069] = 1;
mem[3070] = 1;
mem[3071] = 1;
mem[3072] = 0;
mem[3073] = 0;
mem[3074] = 0;
mem[3075] = 0;
mem[3076] = 0;
mem[3077] = 0;
mem[3078] = 0;
mem[3079] = 0;
mem[3080] = 0;
mem[3081] = 0;
mem[3082] = 0;
mem[3083] = 0;
mem[3084] = 0;
mem[3085] = 0;
mem[3086] = 0;
mem[3087] = 0;
mem[3088] = 0;
mem[3089] = 0;
mem[3090] = 0;
mem[3091] = 0;
mem[3092] = 0;
mem[3093] = 0;
mem[3094] = 0;
mem[3095] = 0;
mem[3096] = 0;
mem[3097] = 0;
mem[3098] = 0;
mem[3099] = 0;
mem[3100] = 0;
mem[3101] = 0;
mem[3102] = 0;
mem[3103] = 0;
mem[3104] = 0;
mem[3105] = 0;
mem[3106] = 0;
mem[3107] = 0;
mem[3108] = 0;
mem[3109] = 0;
mem[3110] = 0;
mem[3111] = 0;
mem[3112] = 0;
mem[3113] = 0;
mem[3114] = 0;
mem[3115] = 0;
mem[3116] = 0;
mem[3117] = 0;
mem[3118] = 0;
mem[3119] = 0;
mem[3120] = 0;
mem[3121] = 0;
mem[3122] = 0;
mem[3123] = 0;
mem[3124] = 0;
mem[3125] = 0;
mem[3126] = 0;
mem[3127] = 0;
mem[3128] = 0;
mem[3129] = 0;
mem[3130] = 0;
mem[3131] = 0;
mem[3132] = 0;
mem[3133] = 0;
mem[3134] = 0;
mem[3135] = 0;
mem[3136] = 0;
mem[3137] = 0;
mem[3138] = 0;
mem[3139] = 0;
mem[3140] = 1;
mem[3141] = 1;
mem[3142] = 1;
mem[3143] = 1;
mem[3144] = 0;
mem[3145] = 0;
mem[3146] = 0;
mem[3147] = 0;
mem[3148] = 0;
mem[3149] = 0;
mem[3150] = 0;
mem[3151] = 0;
mem[3152] = 0;
mem[3153] = 0;
mem[3154] = 0;
mem[3155] = 0;
mem[3156] = 0;
mem[3157] = 0;
mem[3158] = 1;
mem[3159] = 1;
mem[3160] = 1;
mem[3161] = 1;
mem[3162] = 0;
mem[3163] = 0;
mem[3164] = 0;
mem[3165] = 0;
mem[3166] = 0;
mem[3167] = 0;
mem[3168] = 0;
mem[3169] = 0;
mem[3170] = 0;
mem[3171] = 0;
mem[3172] = 0;
mem[3173] = 0;
mem[3174] = 0;
mem[3175] = 0;
mem[3176] = 0;
mem[3177] = 0;
mem[3178] = 0;
mem[3179] = 0;
mem[3180] = 0;
mem[3181] = 0;
mem[3182] = 0;
mem[3183] = 0;
mem[3184] = 0;
mem[3185] = 0;
mem[3186] = 0;
mem[3187] = 0;
mem[3188] = 0;
mem[3189] = 0;
mem[3190] = 0;
mem[3191] = 0;
mem[3192] = 0;
mem[3193] = 0;
mem[3194] = 0;
mem[3195] = 0;
mem[3196] = 0;
mem[3197] = 0;
mem[3198] = 0;
mem[3199] = 0;
mem[3200] = 0;
mem[3201] = 0;
mem[3202] = 0;
mem[3203] = 0;
mem[3204] = 0;
mem[3205] = 0;
mem[3206] = 0;
mem[3207] = 0;
mem[3208] = 0;
mem[3209] = 0;
mem[3210] = 0;
mem[3211] = 0;
mem[3212] = 0;
mem[3213] = 0;
mem[3214] = 0;
mem[3215] = 0;
mem[3216] = 0;
mem[3217] = 0;
mem[3218] = 0;
mem[3219] = 0;
mem[3220] = 0;
mem[3221] = 0;
mem[3222] = 0;
mem[3223] = 0;
mem[3224] = 0;
mem[3225] = 0;
mem[3226] = 0;
mem[3227] = 0;
mem[3228] = 0;
mem[3229] = 0;
mem[3230] = 0;
mem[3231] = 0;
mem[3232] = 1;
mem[3233] = 1;
mem[3234] = 1;
mem[3235] = 0;
mem[3236] = 0;
mem[3237] = 0;
mem[3238] = 0;
mem[3239] = 0;
mem[3240] = 0;
mem[3241] = 0;
mem[3242] = 0;
mem[3243] = 0;
mem[3244] = 0;
mem[3245] = 0;
mem[3246] = 1;
mem[3247] = 1;
mem[3248] = 1;
mem[3249] = 1;
mem[3250] = 1;
mem[3251] = 1;
mem[3252] = 0;
mem[3253] = 0;
mem[3254] = 0;
mem[3255] = 0;
mem[3256] = 0;
mem[3257] = 0;
mem[3258] = 0;
mem[3259] = 0;
mem[3260] = 0;
mem[3261] = 0;
mem[3262] = 0;
mem[3263] = 0;
mem[3264] = 0;
mem[3265] = 0;
mem[3266] = 0;
mem[3267] = 0;
mem[3268] = 0;
mem[3269] = 0;
mem[3270] = 0;
mem[3271] = 0;
mem[3272] = 0;
mem[3273] = 0;
mem[3274] = 0;
mem[3275] = 0;
mem[3276] = 0;
mem[3277] = 0;
mem[3278] = 0;
mem[3279] = 0;
mem[3280] = 0;
mem[3281] = 0;
mem[3282] = 0;
mem[3283] = 0;
mem[3284] = 0;
mem[3285] = 0;
mem[3286] = 0;
mem[3287] = 0;
mem[3288] = 0;
mem[3289] = 0;
mem[3290] = 0;
mem[3291] = 0;
mem[3292] = 0;
mem[3293] = 0;
mem[3294] = 0;
mem[3295] = 0;
mem[3296] = 0;
mem[3297] = 0;
mem[3298] = 0;
mem[3299] = 0;
mem[3300] = 0;
mem[3301] = 0;
mem[3302] = 0;
mem[3303] = 0;
mem[3304] = 0;
mem[3305] = 0;
mem[3306] = 0;
mem[3307] = 0;
mem[3308] = 0;
mem[3309] = 0;
mem[3310] = 0;
mem[3311] = 0;
mem[3312] = 0;
mem[3313] = 0;
mem[3314] = 0;
mem[3315] = 0;
mem[3316] = 0;
mem[3317] = 0;
mem[3318] = 0;
mem[3319] = 0;
mem[3320] = 0;
mem[3321] = 0;
mem[3322] = 0;
mem[3323] = 1;
mem[3324] = 1;
mem[3325] = 1;
mem[3326] = 1;
mem[3327] = 1;
mem[3328] = 0;
mem[3329] = 0;
mem[3330] = 0;
mem[3331] = 0;
mem[3332] = 0;
mem[3333] = 0;
mem[3334] = 0;
mem[3335] = 1;
mem[3336] = 1;
mem[3337] = 1;
mem[3338] = 1;
mem[3339] = 1;
mem[3340] = 0;
mem[3341] = 0;
mem[3342] = 0;
mem[3343] = 0;
mem[3344] = 0;
mem[3345] = 0;
mem[3346] = 0;
mem[3347] = 0;
mem[3348] = 0;
mem[3349] = 0;
mem[3350] = 0;
mem[3351] = 0;
mem[3352] = 0;
mem[3353] = 0;
mem[3354] = 0;
mem[3355] = 0;
mem[3356] = 0;
mem[3357] = 0;
mem[3358] = 0;
mem[3359] = 0;
mem[3360] = 0;
mem[3361] = 0;
mem[3362] = 0;
mem[3363] = 0;
mem[3364] = 0;
mem[3365] = 0;
mem[3366] = 0;
mem[3367] = 0;
mem[3368] = 0;
mem[3369] = 0;
mem[3370] = 0;
mem[3371] = 0;
mem[3372] = 0;
mem[3373] = 0;
mem[3374] = 0;
mem[3375] = 0;
mem[3376] = 0;
mem[3377] = 0;
mem[3378] = 0;
mem[3379] = 0;
mem[3380] = 0;
mem[3381] = 0;
mem[3382] = 0;
mem[3383] = 0;
mem[3384] = 0;
mem[3385] = 0;
mem[3386] = 0;
mem[3387] = 0;
mem[3388] = 0;
mem[3389] = 0;
mem[3390] = 0;
mem[3391] = 0;
mem[3392] = 0;
mem[3393] = 0;
mem[3394] = 0;
mem[3395] = 0;
mem[3396] = 0;
mem[3397] = 0;
mem[3398] = 0;
mem[3399] = 0;
mem[3400] = 0;
mem[3401] = 0;
mem[3402] = 0;
mem[3403] = 0;
mem[3404] = 0;
mem[3405] = 0;
mem[3406] = 0;
mem[3407] = 0;
mem[3408] = 0;
mem[3409] = 0;
mem[3410] = 0;
mem[3411] = 0;
mem[3412] = 0;
mem[3413] = 0;
mem[3414] = 0;
mem[3415] = 1;
mem[3416] = 1;
mem[3417] = 1;
mem[3418] = 0;
mem[3419] = 0;
mem[3420] = 0;
mem[3421] = 0;
mem[3422] = 0;
mem[3423] = 1;
mem[3424] = 1;
mem[3425] = 1;
mem[3426] = 1;
mem[3427] = 1;
mem[3428] = 0;
mem[3429] = 0;
mem[3430] = 0;
mem[3431] = 0;
mem[3432] = 0;
mem[3433] = 0;
mem[3434] = 0;
mem[3435] = 0;
mem[3436] = 0;
mem[3437] = 0;
mem[3438] = 0;
mem[3439] = 0;
mem[3440] = 0;
mem[3441] = 0;
mem[3442] = 0;
mem[3443] = 0;
mem[3444] = 0;
mem[3445] = 0;
mem[3446] = 0;
mem[3447] = 0;
mem[3448] = 0;
mem[3449] = 0;
mem[3450] = 0;
mem[3451] = 0;
mem[3452] = 0;
mem[3453] = 0;
mem[3454] = 0;
mem[3455] = 0;
mem[3456] = 0;
mem[3457] = 0;
mem[3458] = 0;
mem[3459] = 0;
mem[3460] = 0;
mem[3461] = 0;
mem[3462] = 0;
mem[3463] = 0;
mem[3464] = 0;
mem[3465] = 0;
mem[3466] = 0;
mem[3467] = 0;
mem[3468] = 0;
mem[3469] = 0;
mem[3470] = 0;
mem[3471] = 0;
mem[3472] = 0;
mem[3473] = 0;
mem[3474] = 0;
mem[3475] = 0;
mem[3476] = 0;
mem[3477] = 0;
mem[3478] = 0;
mem[3479] = 0;
mem[3480] = 0;
mem[3481] = 0;
mem[3482] = 0;
mem[3483] = 0;
mem[3484] = 0;
mem[3485] = 0;
mem[3486] = 0;
mem[3487] = 0;
mem[3488] = 0;
mem[3489] = 0;
mem[3490] = 0;
mem[3491] = 0;
mem[3492] = 0;
mem[3493] = 0;
mem[3494] = 0;
mem[3495] = 0;
mem[3496] = 0;
mem[3497] = 0;
mem[3498] = 0;
mem[3499] = 0;
mem[3500] = 0;
mem[3501] = 1;
mem[3502] = 1;
mem[3503] = 1;
mem[3504] = 1;
mem[3505] = 1;
mem[3506] = 1;
mem[3507] = 1;
mem[3508] = 0;
mem[3509] = 0;
mem[3510] = 0;
mem[3511] = 1;
mem[3512] = 1;
mem[3513] = 1;
mem[3514] = 1;
mem[3515] = 1;
mem[3516] = 0;
mem[3517] = 0;
mem[3518] = 0;
mem[3519] = 0;
mem[3520] = 0;
mem[3521] = 0;
mem[3522] = 0;
mem[3523] = 0;
mem[3524] = 0;
mem[3525] = 0;
mem[3526] = 0;
mem[3527] = 0;
mem[3528] = 0;
mem[3529] = 0;
mem[3530] = 0;
mem[3531] = 0;
mem[3532] = 0;
mem[3533] = 0;
mem[3534] = 0;
mem[3535] = 0;
mem[3536] = 0;
mem[3537] = 0;
mem[3538] = 0;
mem[3539] = 0;
mem[3540] = 0;
mem[3541] = 0;
mem[3542] = 0;
mem[3543] = 0;
mem[3544] = 0;
mem[3545] = 0;
mem[3546] = 0;
mem[3547] = 0;
mem[3548] = 0;
mem[3549] = 0;
mem[3550] = 0;
mem[3551] = 0;
mem[3552] = 0;
mem[3553] = 0;
mem[3554] = 0;
mem[3555] = 0;
mem[3556] = 0;
mem[3557] = 0;
mem[3558] = 0;
mem[3559] = 0;
mem[3560] = 0;
mem[3561] = 0;
mem[3562] = 0;
mem[3563] = 0;
mem[3564] = 0;
mem[3565] = 0;
mem[3566] = 0;
mem[3567] = 0;
mem[3568] = 0;
mem[3569] = 0;
mem[3570] = 0;
mem[3571] = 0;
mem[3572] = 0;
mem[3573] = 0;
mem[3574] = 0;
mem[3575] = 0;
mem[3576] = 0;
mem[3577] = 0;
mem[3578] = 0;
mem[3579] = 0;
mem[3580] = 0;
mem[3581] = 0;
mem[3582] = 0;
mem[3583] = 0;
mem[3584] = 0;
mem[3585] = 0;
mem[3586] = 0;
mem[3587] = 0;
mem[3588] = 0;
mem[3589] = 1;
mem[3590] = 1;
mem[3591] = 1;
mem[3592] = 1;
mem[3593] = 1;
mem[3594] = 1;
mem[3595] = 1;
mem[3596] = 0;
mem[3597] = 0;
mem[3598] = 0;
mem[3599] = 0;
mem[3600] = 0;
mem[3601] = 1;
mem[3602] = 1;
mem[3603] = 1;
mem[3604] = 1;
mem[3605] = 1;
mem[3606] = 0;
mem[3607] = 0;
mem[3608] = 0;
mem[3609] = 0;
mem[3610] = 0;
mem[3611] = 0;
mem[3612] = 0;
mem[3613] = 0;
mem[3614] = 0;
mem[3615] = 0;
mem[3616] = 0;
mem[3617] = 0;
mem[3618] = 0;
mem[3619] = 0;
mem[3620] = 0;
mem[3621] = 0;
mem[3622] = 0;
mem[3623] = 0;
mem[3624] = 0;
mem[3625] = 0;
mem[3626] = 0;
mem[3627] = 0;
mem[3628] = 0;
mem[3629] = 0;
mem[3630] = 0;
mem[3631] = 0;
mem[3632] = 0;
mem[3633] = 0;
mem[3634] = 0;
mem[3635] = 0;
mem[3636] = 0;
mem[3637] = 0;
mem[3638] = 0;
mem[3639] = 0;
mem[3640] = 0;
mem[3641] = 0;
mem[3642] = 0;
mem[3643] = 0;
mem[3644] = 0;
mem[3645] = 0;
mem[3646] = 0;
mem[3647] = 0;
mem[3648] = 0;
mem[3649] = 0;
mem[3650] = 0;
mem[3651] = 0;
mem[3652] = 0;
mem[3653] = 0;
mem[3654] = 0;
mem[3655] = 0;
mem[3656] = 0;
mem[3657] = 0;
mem[3658] = 0;
mem[3659] = 0;
mem[3660] = 0;
mem[3661] = 0;
mem[3662] = 0;
mem[3663] = 0;
mem[3664] = 0;
mem[3665] = 0;
mem[3666] = 0;
mem[3667] = 0;
mem[3668] = 0;
mem[3669] = 0;
mem[3670] = 0;
mem[3671] = 0;
mem[3672] = 0;
mem[3673] = 0;
mem[3674] = 0;
mem[3675] = 0;
mem[3676] = 0;
mem[3677] = 0;
mem[3678] = 0;
mem[3679] = 1;
mem[3680] = 1;
mem[3681] = 1;
mem[3682] = 1;
mem[3683] = 1;
mem[3684] = 1;
mem[3685] = 0;
mem[3686] = 0;
mem[3687] = 0;
mem[3688] = 0;
mem[3689] = 0;
mem[3690] = 0;
mem[3691] = 1;
mem[3692] = 1;
mem[3693] = 1;
mem[3694] = 1;
mem[3695] = 1;
mem[3696] = 1;
mem[3697] = 1;
mem[3698] = 1;
mem[3699] = 1;
mem[3700] = 1;
mem[3701] = 1;
mem[3702] = 1;
mem[3703] = 0;
mem[3704] = 0;
mem[3705] = 0;
mem[3706] = 0;
mem[3707] = 0;
mem[3708] = 0;
mem[3709] = 0;
mem[3710] = 0;
mem[3711] = 0;
mem[3712] = 0;
mem[3713] = 0;
mem[3714] = 0;
mem[3715] = 0;
mem[3716] = 0;
mem[3717] = 0;
mem[3718] = 0;
mem[3719] = 0;
mem[3720] = 0;
mem[3721] = 0;
mem[3722] = 0;
mem[3723] = 0;
mem[3724] = 0;
mem[3725] = 0;
mem[3726] = 0;
mem[3727] = 0;
mem[3728] = 0;
mem[3729] = 0;
mem[3730] = 0;
mem[3731] = 0;
mem[3732] = 0;
mem[3733] = 0;
mem[3734] = 0;
mem[3735] = 0;
mem[3736] = 0;
mem[3737] = 0;
mem[3738] = 0;
mem[3739] = 0;
mem[3740] = 0;
mem[3741] = 0;
mem[3742] = 0;
mem[3743] = 0;
mem[3744] = 0;
mem[3745] = 0;
mem[3746] = 0;
mem[3747] = 0;
mem[3748] = 0;
mem[3749] = 0;
mem[3750] = 0;
mem[3751] = 0;
mem[3752] = 0;
mem[3753] = 0;
mem[3754] = 0;
mem[3755] = 0;
mem[3756] = 0;
mem[3757] = 0;
mem[3758] = 0;
mem[3759] = 0;
mem[3760] = 0;
mem[3761] = 0;
mem[3762] = 0;
mem[3763] = 0;
mem[3764] = 0;
mem[3765] = 0;
mem[3766] = 0;
mem[3767] = 0;
mem[3768] = 1;
mem[3769] = 1;
mem[3770] = 1;
mem[3771] = 0;
mem[3772] = 0;
mem[3773] = 0;
mem[3774] = 0;
mem[3775] = 0;
mem[3776] = 0;
mem[3777] = 0;
mem[3778] = 0;
mem[3779] = 0;
mem[3780] = 0;
mem[3781] = 0;
mem[3782] = 0;
mem[3783] = 0;
mem[3784] = 0;
mem[3785] = 0;
mem[3786] = 1;
mem[3787] = 1;
mem[3788] = 1;
mem[3789] = 1;
mem[3790] = 1;
mem[3791] = 1;
mem[3792] = 1;
mem[3793] = 0;
mem[3794] = 0;
mem[3795] = 0;
mem[3796] = 0;
mem[3797] = 0;
mem[3798] = 0;
mem[3799] = 0;
mem[3800] = 0;
mem[3801] = 0;
mem[3802] = 0;
mem[3803] = 0;
mem[3804] = 0;
mem[3805] = 0;
mem[3806] = 0;
mem[3807] = 0;
mem[3808] = 0;
mem[3809] = 0;
mem[3810] = 0;
mem[3811] = 0;
mem[3812] = 0;
mem[3813] = 0;
mem[3814] = 0;
mem[3815] = 0;
mem[3816] = 0;
mem[3817] = 0;
mem[3818] = 0;
mem[3819] = 0;
mem[3820] = 0;
mem[3821] = 0;
mem[3822] = 0;
mem[3823] = 0;
mem[3824] = 0;
mem[3825] = 0;
mem[3826] = 0;
mem[3827] = 0;
mem[3828] = 0;
mem[3829] = 0;
mem[3830] = 0;
mem[3831] = 0;
mem[3832] = 0;
mem[3833] = 0;
mem[3834] = 0;
mem[3835] = 0;
mem[3836] = 1;
mem[3837] = 1;
mem[3838] = 0;
mem[3839] = 0;
mem[3840] = 0;
mem[3841] = 0;
mem[3842] = 0;
mem[3843] = 0;
mem[3844] = 1;
mem[3845] = 1;
mem[3846] = 1;
mem[3847] = 0;
mem[3848] = 0;
mem[3849] = 0;
mem[3850] = 0;
mem[3851] = 0;
mem[3852] = 0;
mem[3853] = 1;
mem[3854] = 1;
mem[3855] = 0;
mem[3856] = 0;
mem[3857] = 0;
mem[3858] = 1;
mem[3859] = 1;
mem[3860] = 1;
mem[3861] = 0;
mem[3862] = 0;
mem[3863] = 0;
mem[3864] = 0;
mem[3865] = 0;
mem[3866] = 0;
mem[3867] = 0;
mem[3868] = 0;
mem[3869] = 0;
mem[3870] = 0;
mem[3871] = 0;
mem[3872] = 0;
mem[3873] = 0;
mem[3874] = 0;
mem[3875] = 0;
mem[3876] = 0;
mem[3877] = 0;
mem[3878] = 0;
mem[3879] = 0;
mem[3880] = 1;
mem[3881] = 1;
mem[3882] = 1;
mem[3883] = 0;
mem[3884] = 0;
mem[3885] = 0;
mem[3886] = 0;
mem[3887] = 0;
mem[3888] = 0;
mem[3889] = 0;
mem[3890] = 0;
mem[3891] = 0;
mem[3892] = 0;
mem[3893] = 0;
mem[3894] = 0;
mem[3895] = 0;
mem[3896] = 0;
mem[3897] = 0;
mem[3898] = 0;
mem[3899] = 0;
mem[3900] = 0;
mem[3901] = 0;
mem[3902] = 0;
mem[3903] = 0;
mem[3904] = 0;
mem[3905] = 0;
mem[3906] = 0;
mem[3907] = 1;
mem[3908] = 1;
mem[3909] = 1;
mem[3910] = 0;
mem[3911] = 0;
mem[3912] = 0;
mem[3913] = 0;
mem[3914] = 0;
mem[3915] = 0;
mem[3916] = 0;
mem[3917] = 1;
mem[3918] = 0;
mem[3919] = 0;
mem[3920] = 0;
mem[3921] = 0;
mem[3922] = 0;
mem[3923] = 0;
mem[3924] = 0;
mem[3925] = 1;
mem[3926] = 1;
mem[3927] = 1;
mem[3928] = 1;
mem[3929] = 0;
mem[3930] = 0;
mem[3931] = 0;
mem[3932] = 0;
mem[3933] = 0;
mem[3934] = 1;
mem[3935] = 1;
mem[3936] = 1;
mem[3937] = 0;
mem[3938] = 0;
mem[3939] = 0;
mem[3940] = 0;
mem[3941] = 0;
mem[3942] = 1;
mem[3943] = 1;
mem[3944] = 1;
mem[3945] = 1;
mem[3946] = 0;
mem[3947] = 0;
mem[3948] = 0;
mem[3949] = 0;
mem[3950] = 1;
mem[3951] = 1;
mem[3952] = 0;
mem[3953] = 0;
mem[3954] = 0;
mem[3955] = 0;
mem[3956] = 0;
mem[3957] = 0;
mem[3958] = 0;
mem[3959] = 0;
mem[3960] = 0;
mem[3961] = 0;
mem[3962] = 0;
mem[3963] = 0;
mem[3964] = 0;
mem[3965] = 0;
mem[3966] = 0;
mem[3967] = 0;
mem[3968] = 0;
mem[3969] = 1;
mem[3970] = 1;
mem[3971] = 1;
mem[3972] = 0;
mem[3973] = 0;
mem[3974] = 0;
mem[3975] = 0;
mem[3976] = 0;
mem[3977] = 0;
mem[3978] = 0;
mem[3979] = 0;
mem[3980] = 0;
mem[3981] = 0;
mem[3982] = 0;
mem[3983] = 0;
mem[3984] = 0;
mem[3985] = 0;
mem[3986] = 0;
mem[3987] = 0;
mem[3988] = 0;
mem[3989] = 0;
mem[3990] = 0;
mem[3991] = 0;
mem[3992] = 0;
mem[3993] = 0;
mem[3994] = 0;
mem[3995] = 0;
mem[3996] = 0;
mem[3997] = 1;
mem[3998] = 1;
mem[3999] = 1;
mem[4000] = 0;
mem[4001] = 0;
mem[4002] = 0;
mem[4003] = 0;
mem[4004] = 0;
mem[4005] = 0;
mem[4006] = 1;
mem[4007] = 1;
mem[4008] = 1;
mem[4009] = 0;
mem[4010] = 0;
mem[4011] = 0;
mem[4012] = 0;
mem[4013] = 0;
mem[4014] = 0;
mem[4015] = 1;
mem[4016] = 1;
mem[4017] = 1;
mem[4018] = 1;
mem[4019] = 1;
mem[4020] = 0;
mem[4021] = 0;
mem[4022] = 0;
mem[4023] = 0;
mem[4024] = 1;
mem[4025] = 1;
mem[4026] = 1;
mem[4027] = 1;
mem[4028] = 0;
mem[4029] = 0;
mem[4030] = 0;
mem[4031] = 0;
mem[4032] = 1;
mem[4033] = 1;
mem[4034] = 1;
mem[4035] = 1;
mem[4036] = 1;
mem[4037] = 0;
mem[4038] = 0;
mem[4039] = 0;
mem[4040] = 1;
mem[4041] = 1;
mem[4042] = 0;
mem[4043] = 0;
mem[4044] = 0;
mem[4045] = 0;
mem[4046] = 0;
mem[4047] = 0;
mem[4048] = 0;
mem[4049] = 0;
mem[4050] = 0;
mem[4051] = 0;
mem[4052] = 0;
mem[4053] = 0;
mem[4054] = 0;
mem[4055] = 0;
mem[4056] = 0;
mem[4057] = 0;
mem[4058] = 0;
mem[4059] = 1;
mem[4060] = 1;
mem[4061] = 1;
mem[4062] = 0;
mem[4063] = 0;
mem[4064] = 0;
mem[4065] = 0;
mem[4066] = 0;
mem[4067] = 0;
mem[4068] = 0;
mem[4069] = 0;
mem[4070] = 0;
mem[4071] = 0;
mem[4072] = 1;
mem[4073] = 1;
mem[4074] = 1;
mem[4075] = 0;
mem[4076] = 0;
mem[4077] = 0;
mem[4078] = 0;
mem[4079] = 1;
mem[4080] = 1;
mem[4081] = 1;
mem[4082] = 0;
mem[4083] = 0;
mem[4084] = 0;
mem[4085] = 0;
mem[4086] = 0;
mem[4087] = 1;
mem[4088] = 1;
mem[4089] = 1;
mem[4090] = 0;
mem[4091] = 0;
mem[4092] = 0;
mem[4093] = 0;
mem[4094] = 0;
mem[4095] = 1;
mem[4096] = 1;
mem[4097] = 1;
mem[4098] = 1;
mem[4099] = 0;
mem[4100] = 0;
mem[4101] = 0;
mem[4102] = 0;
mem[4103] = 0;
mem[4104] = 0;
mem[4105] = 1;
mem[4106] = 1;
mem[4107] = 1;
mem[4108] = 1;
mem[4109] = 1;
mem[4110] = 0;
mem[4111] = 0;
mem[4112] = 0;
mem[4113] = 1;
mem[4114] = 1;
mem[4115] = 1;
mem[4116] = 1;
mem[4117] = 1;
mem[4118] = 0;
mem[4119] = 0;
mem[4120] = 0;
mem[4121] = 0;
mem[4122] = 1;
mem[4123] = 1;
mem[4124] = 0;
mem[4125] = 1;
mem[4126] = 1;
mem[4127] = 1;
mem[4128] = 1;
mem[4129] = 0;
mem[4130] = 1;
mem[4131] = 1;
mem[4132] = 0;
mem[4133] = 0;
mem[4134] = 0;
mem[4135] = 0;
mem[4136] = 0;
mem[4137] = 0;
mem[4138] = 0;
mem[4139] = 0;
mem[4140] = 0;
mem[4141] = 0;
mem[4142] = 0;
mem[4143] = 0;
mem[4144] = 0;
mem[4145] = 0;
mem[4146] = 0;
mem[4147] = 0;
mem[4148] = 0;
mem[4149] = 1;
mem[4150] = 1;
mem[4151] = 1;
mem[4152] = 0;
mem[4153] = 1;
mem[4154] = 1;
mem[4155] = 1;
mem[4156] = 0;
mem[4157] = 0;
mem[4158] = 0;
mem[4159] = 0;
mem[4160] = 0;
mem[4161] = 1;
mem[4162] = 1;
mem[4163] = 1;
mem[4164] = 1;
mem[4165] = 0;
mem[4166] = 0;
mem[4167] = 0;
mem[4168] = 0;
mem[4169] = 1;
mem[4170] = 1;
mem[4171] = 1;
mem[4172] = 1;
mem[4173] = 0;
mem[4174] = 0;
mem[4175] = 0;
mem[4176] = 0;
mem[4177] = 1;
mem[4178] = 1;
mem[4179] = 1;
mem[4180] = 1;
mem[4181] = 1;
mem[4182] = 0;
mem[4183] = 0;
mem[4184] = 0;
mem[4185] = 1;
mem[4186] = 1;
mem[4187] = 1;
mem[4188] = 1;
mem[4189] = 1;
mem[4190] = 0;
mem[4191] = 0;
mem[4192] = 0;
mem[4193] = 0;
mem[4194] = 1;
mem[4195] = 1;
mem[4196] = 0;
mem[4197] = 1;
mem[4198] = 1;
mem[4199] = 1;
mem[4200] = 0;
mem[4201] = 0;
mem[4202] = 0;
mem[4203] = 1;
mem[4204] = 1;
mem[4205] = 0;
mem[4206] = 0;
mem[4207] = 1;
mem[4208] = 1;
mem[4209] = 0;
mem[4210] = 0;
mem[4211] = 1;
mem[4212] = 1;
mem[4213] = 0;
mem[4214] = 0;
mem[4215] = 0;
mem[4216] = 0;
mem[4217] = 1;
mem[4218] = 1;
mem[4219] = 1;
mem[4220] = 1;
mem[4221] = 1;
mem[4222] = 1;
mem[4223] = 0;
mem[4224] = 0;
mem[4225] = 0;
mem[4226] = 0;
mem[4227] = 0;
mem[4228] = 0;
mem[4229] = 0;
mem[4230] = 0;
mem[4231] = 0;
mem[4232] = 0;
mem[4233] = 0;
mem[4234] = 0;
mem[4235] = 0;
mem[4236] = 0;
mem[4237] = 0;
mem[4238] = 1;
mem[4239] = 1;
mem[4240] = 1;
mem[4241] = 0;
mem[4242] = 1;
mem[4243] = 1;
mem[4244] = 1;
mem[4245] = 1;
mem[4246] = 0;
mem[4247] = 0;
mem[4248] = 0;
mem[4249] = 0;
mem[4250] = 0;
mem[4251] = 1;
mem[4252] = 1;
mem[4253] = 1;
mem[4254] = 1;
mem[4255] = 1;
mem[4256] = 0;
mem[4257] = 0;
mem[4258] = 1;
mem[4259] = 1;
mem[4260] = 1;
mem[4261] = 1;
mem[4262] = 1;
mem[4263] = 0;
mem[4264] = 0;
mem[4265] = 0;
mem[4266] = 1;
mem[4267] = 1;
mem[4268] = 0;
mem[4269] = 1;
mem[4270] = 1;
mem[4271] = 1;
mem[4272] = 0;
mem[4273] = 0;
mem[4274] = 1;
mem[4275] = 1;
mem[4276] = 1;
mem[4277] = 0;
mem[4278] = 1;
mem[4279] = 1;
mem[4280] = 1;
mem[4281] = 0;
mem[4282] = 0;
mem[4283] = 0;
mem[4284] = 1;
mem[4285] = 1;
mem[4286] = 0;
mem[4287] = 0;
mem[4288] = 1;
mem[4289] = 1;
mem[4290] = 1;
mem[4291] = 0;
mem[4292] = 1;
mem[4293] = 1;
mem[4294] = 1;
mem[4295] = 0;
mem[4296] = 0;
mem[4297] = 1;
mem[4298] = 1;
mem[4299] = 0;
mem[4300] = 1;
mem[4301] = 1;
mem[4302] = 0;
mem[4303] = 0;
mem[4304] = 0;
mem[4305] = 0;
mem[4306] = 0;
mem[4307] = 0;
mem[4308] = 1;
mem[4309] = 1;
mem[4310] = 1;
mem[4311] = 1;
mem[4312] = 1;
mem[4313] = 0;
mem[4314] = 0;
mem[4315] = 0;
mem[4316] = 0;
mem[4317] = 0;
mem[4318] = 0;
mem[4319] = 0;
mem[4320] = 0;
mem[4321] = 0;
mem[4322] = 0;
mem[4323] = 0;
mem[4324] = 0;
mem[4325] = 0;
mem[4326] = 0;
mem[4327] = 0;
mem[4328] = 1;
mem[4329] = 1;
mem[4330] = 0;
mem[4331] = 1;
mem[4332] = 1;
mem[4333] = 1;
mem[4334] = 1;
mem[4335] = 1;
mem[4336] = 1;
mem[4337] = 0;
mem[4338] = 0;
mem[4339] = 0;
mem[4340] = 1;
mem[4341] = 1;
mem[4342] = 1;
mem[4343] = 1;
mem[4344] = 1;
mem[4345] = 1;
mem[4346] = 0;
mem[4347] = 0;
mem[4348] = 1;
mem[4349] = 1;
mem[4350] = 1;
mem[4351] = 1;
mem[4352] = 1;
mem[4353] = 1;
mem[4354] = 0;
mem[4355] = 1;
mem[4356] = 1;
mem[4357] = 0;
mem[4358] = 0;
mem[4359] = 1;
mem[4360] = 1;
mem[4361] = 1;
mem[4362] = 1;
mem[4363] = 0;
mem[4364] = 1;
mem[4365] = 1;
mem[4366] = 0;
mem[4367] = 0;
mem[4368] = 0;
mem[4369] = 1;
mem[4370] = 1;
mem[4371] = 0;
mem[4372] = 1;
mem[4373] = 1;
mem[4374] = 1;
mem[4375] = 0;
mem[4376] = 0;
mem[4377] = 0;
mem[4378] = 1;
mem[4379] = 1;
mem[4380] = 1;
mem[4381] = 0;
mem[4382] = 1;
mem[4383] = 1;
mem[4384] = 0;
mem[4385] = 0;
mem[4386] = 0;
mem[4387] = 1;
mem[4388] = 1;
mem[4389] = 1;
mem[4390] = 1;
mem[4391] = 0;
mem[4392] = 0;
mem[4393] = 0;
mem[4394] = 0;
mem[4395] = 0;
mem[4396] = 0;
mem[4397] = 0;
mem[4398] = 0;
mem[4399] = 0;
mem[4400] = 1;
mem[4401] = 1;
mem[4402] = 1;
mem[4403] = 0;
mem[4404] = 0;
mem[4405] = 0;
mem[4406] = 0;
mem[4407] = 0;
mem[4408] = 0;
mem[4409] = 0;
mem[4410] = 0;
mem[4411] = 0;
mem[4412] = 0;
mem[4413] = 0;
mem[4414] = 0;
mem[4415] = 0;
mem[4416] = 0;
mem[4417] = 0;
mem[4418] = 1;
mem[4419] = 1;
mem[4420] = 1;
mem[4421] = 1;
mem[4422] = 1;
mem[4423] = 1;
mem[4424] = 0;
mem[4425] = 1;
mem[4426] = 1;
mem[4427] = 0;
mem[4428] = 0;
mem[4429] = 0;
mem[4430] = 1;
mem[4431] = 1;
mem[4432] = 0;
mem[4433] = 0;
mem[4434] = 1;
mem[4435] = 1;
mem[4436] = 1;
mem[4437] = 0;
mem[4438] = 1;
mem[4439] = 1;
mem[4440] = 0;
mem[4441] = 0;
mem[4442] = 1;
mem[4443] = 1;
mem[4444] = 0;
mem[4445] = 1;
mem[4446] = 1;
mem[4447] = 0;
mem[4448] = 0;
mem[4449] = 0;
mem[4450] = 1;
mem[4451] = 1;
mem[4452] = 1;
mem[4453] = 1;
mem[4454] = 1;
mem[4455] = 1;
mem[4456] = 0;
mem[4457] = 0;
mem[4458] = 0;
mem[4459] = 1;
mem[4460] = 1;
mem[4461] = 1;
mem[4462] = 1;
mem[4463] = 1;
mem[4464] = 0;
mem[4465] = 0;
mem[4466] = 0;
mem[4467] = 0;
mem[4468] = 1;
mem[4469] = 1;
mem[4470] = 1;
mem[4471] = 1;
mem[4472] = 1;
mem[4473] = 1;
mem[4474] = 0;
mem[4475] = 0;
mem[4476] = 0;
mem[4477] = 0;
mem[4478] = 1;
mem[4479] = 1;
mem[4480] = 1;
mem[4481] = 0;
mem[4482] = 0;
mem[4483] = 0;
mem[4484] = 0;
mem[4485] = 0;
mem[4486] = 0;
mem[4487] = 0;
mem[4488] = 0;
mem[4489] = 0;
mem[4490] = 0;
mem[4491] = 0;
mem[4492] = 0;
mem[4493] = 0;
mem[4494] = 0;
mem[4495] = 0;
mem[4496] = 0;
mem[4497] = 0;
mem[4498] = 0;
mem[4499] = 0;
mem[4500] = 0;
mem[4501] = 0;
mem[4502] = 0;
mem[4503] = 0;
mem[4504] = 0;
mem[4505] = 0;
mem[4506] = 0;
mem[4507] = 0;
mem[4508] = 1;
mem[4509] = 1;
mem[4510] = 1;
mem[4511] = 1;
mem[4512] = 0;
mem[4513] = 0;
mem[4514] = 0;
mem[4515] = 1;
mem[4516] = 1;
mem[4517] = 1;
mem[4518] = 0;
mem[4519] = 1;
mem[4520] = 1;
mem[4521] = 1;
mem[4522] = 0;
mem[4523] = 0;
mem[4524] = 1;
mem[4525] = 1;
mem[4526] = 1;
mem[4527] = 1;
mem[4528] = 1;
mem[4529] = 1;
mem[4530] = 0;
mem[4531] = 0;
mem[4532] = 1;
mem[4533] = 1;
mem[4534] = 1;
mem[4535] = 0;
mem[4536] = 1;
mem[4537] = 0;
mem[4538] = 0;
mem[4539] = 0;
mem[4540] = 1;
mem[4541] = 1;
mem[4542] = 1;
mem[4543] = 1;
mem[4544] = 1;
mem[4545] = 0;
mem[4546] = 0;
mem[4547] = 0;
mem[4548] = 0;
mem[4549] = 0;
mem[4550] = 1;
mem[4551] = 1;
mem[4552] = 1;
mem[4553] = 1;
mem[4554] = 0;
mem[4555] = 0;
mem[4556] = 0;
mem[4557] = 0;
mem[4558] = 1;
mem[4559] = 1;
mem[4560] = 1;
mem[4561] = 1;
mem[4562] = 1;
mem[4563] = 0;
mem[4564] = 0;
mem[4565] = 0;
mem[4566] = 0;
mem[4567] = 0;
mem[4568] = 1;
mem[4569] = 1;
mem[4570] = 0;
mem[4571] = 0;
mem[4572] = 0;
mem[4573] = 0;
mem[4574] = 0;
mem[4575] = 0;
mem[4576] = 0;
mem[4577] = 0;
mem[4578] = 0;
mem[4579] = 0;
mem[4580] = 0;
mem[4581] = 0;
mem[4582] = 0;
mem[4583] = 0;
mem[4584] = 0;
mem[4585] = 0;
mem[4586] = 0;
mem[4587] = 0;
mem[4588] = 0;
mem[4589] = 0;
mem[4590] = 0;
mem[4591] = 0;
mem[4592] = 0;
mem[4593] = 0;
mem[4594] = 0;
mem[4595] = 0;
mem[4596] = 0;
mem[4597] = 1;
mem[4598] = 1;
mem[4599] = 1;
mem[4600] = 1;
mem[4601] = 1;
mem[4602] = 0;
mem[4603] = 0;
mem[4604] = 0;
mem[4605] = 0;
mem[4606] = 1;
mem[4607] = 1;
mem[4608] = 1;
mem[4609] = 1;
mem[4610] = 1;
mem[4611] = 0;
mem[4612] = 0;
mem[4613] = 0;
mem[4614] = 0;
mem[4615] = 1;
mem[4616] = 1;
mem[4617] = 1;
mem[4618] = 1;
mem[4619] = 1;
mem[4620] = 0;
mem[4621] = 0;
mem[4622] = 0;
mem[4623] = 1;
mem[4624] = 1;
mem[4625] = 1;
mem[4626] = 1;
mem[4627] = 0;
mem[4628] = 0;
mem[4629] = 0;
mem[4630] = 0;
mem[4631] = 1;
mem[4632] = 1;
mem[4633] = 1;
mem[4634] = 1;
mem[4635] = 0;
mem[4636] = 0;
mem[4637] = 0;
mem[4638] = 0;
mem[4639] = 0;
mem[4640] = 1;
mem[4641] = 1;
mem[4642] = 1;
mem[4643] = 1;
mem[4644] = 0;
mem[4645] = 0;
mem[4646] = 0;
mem[4647] = 0;
mem[4648] = 0;
mem[4649] = 1;
mem[4650] = 1;
mem[4651] = 1;
mem[4652] = 1;
mem[4653] = 0;
mem[4654] = 0;
mem[4655] = 0;
mem[4656] = 0;
mem[4657] = 0;
mem[4658] = 0;
mem[4659] = 0;
mem[4660] = 0;
mem[4661] = 0;
mem[4662] = 0;
mem[4663] = 0;
mem[4664] = 0;
mem[4665] = 0;
mem[4666] = 0;
mem[4667] = 0;
mem[4668] = 0;
mem[4669] = 0;
mem[4670] = 0;
mem[4671] = 0;
mem[4672] = 0;
mem[4673] = 0;
mem[4674] = 0;
mem[4675] = 0;
mem[4676] = 0;
mem[4677] = 0;
mem[4678] = 0;
mem[4679] = 0;
mem[4680] = 0;
mem[4681] = 0;
mem[4682] = 0;
mem[4683] = 0;
mem[4684] = 0;
mem[4685] = 0;
mem[4686] = 0;
mem[4687] = 1;
mem[4688] = 1;
mem[4689] = 1;
mem[4690] = 1;
mem[4691] = 0;
mem[4692] = 0;
mem[4693] = 0;
mem[4694] = 0;
mem[4695] = 0;
mem[4696] = 1;
mem[4697] = 1;
mem[4698] = 1;
mem[4699] = 1;
mem[4700] = 0;
mem[4701] = 0;
mem[4702] = 0;
mem[4703] = 0;
mem[4704] = 0;
mem[4705] = 1;
mem[4706] = 1;
mem[4707] = 1;
mem[4708] = 1;
mem[4709] = 0;
mem[4710] = 0;
mem[4711] = 0;
mem[4712] = 0;
mem[4713] = 1;
mem[4714] = 1;
mem[4715] = 1;
mem[4716] = 1;
mem[4717] = 0;
mem[4718] = 0;
mem[4719] = 0;
mem[4720] = 0;
mem[4721] = 0;
mem[4722] = 1;
mem[4723] = 1;
mem[4724] = 0;
mem[4725] = 0;
mem[4726] = 0;
mem[4727] = 0;
mem[4728] = 0;
mem[4729] = 0;
mem[4730] = 0;
mem[4731] = 1;
mem[4732] = 1;
mem[4733] = 0;
mem[4734] = 0;
mem[4735] = 0;
mem[4736] = 0;
mem[4737] = 0;
mem[4738] = 0;
mem[4739] = 0;
mem[4740] = 1;
mem[4741] = 1;
mem[4742] = 0;
mem[4743] = 0;
mem[4744] = 0;
mem[4745] = 0;
mem[4746] = 0;
mem[4747] = 0;
mem[4748] = 0;
mem[4749] = 0;
mem[4750] = 0;
mem[4751] = 0;
mem[4752] = 0;
mem[4753] = 0;
mem[4754] = 0;
mem[4755] = 0;
mem[4756] = 0;
mem[4757] = 0;
mem[4758] = 0;
mem[4759] = 0;
mem[4760] = 0;
mem[4761] = 0;
mem[4762] = 0;
mem[4763] = 0;
mem[4764] = 0;
mem[4765] = 0;
mem[4766] = 0;
mem[4767] = 0;
mem[4768] = 0;
mem[4769] = 0;
mem[4770] = 0;
mem[4771] = 0;
mem[4772] = 0;
mem[4773] = 0;
mem[4774] = 0;
mem[4775] = 0;
mem[4776] = 0;
mem[4777] = 1;
mem[4778] = 1;
mem[4779] = 0;
mem[4780] = 0;
mem[4781] = 0;
mem[4782] = 0;
mem[4783] = 0;
mem[4784] = 0;
mem[4785] = 0;
mem[4786] = 0;
mem[4787] = 1;
mem[4788] = 1;
mem[4789] = 0;
mem[4790] = 0;
mem[4791] = 0;
mem[4792] = 0;
mem[4793] = 0;
mem[4794] = 0;
mem[4795] = 0;
mem[4796] = 1;
mem[4797] = 1;
mem[4798] = 1;
mem[4799] = 0;
mem[4800] = 0;
mem[4801] = 0;
mem[4802] = 0;
mem[4803] = 0;
mem[4804] = 1;
mem[4805] = 1;
mem[4806] = 0;
mem[4807] = 0;
mem[4808] = 0;
mem[4809] = 0;
mem[4810] = 0;
mem[4811] = 0;
mem[4812] = 1;
mem[4813] = 0;
mem[4814] = 0;
mem[4815] = 0;
mem[4816] = 0;
mem[4817] = 0;
mem[4818] = 0;
mem[4819] = 0;
mem[4820] = 0;
mem[4821] = 0;
mem[4822] = 1;
mem[4823] = 0;
mem[4824] = 0;
mem[4825] = 0;
mem[4826] = 0;
mem[4827] = 0;
mem[4828] = 0;
mem[4829] = 0;
mem[4830] = 1;
mem[4831] = 1;
mem[4832] = 0;
mem[4833] = 0;
mem[4834] = 0;
mem[4835] = 0;
mem[4836] = 0;
mem[4837] = 0;
mem[4838] = 0;
mem[4839] = 0;
mem[4840] = 0;
mem[4841] = 0;
mem[4842] = 0;
mem[4843] = 0;
mem[4844] = 0;
mem[4845] = 0;
mem[4846] = 0;
mem[4847] = 0;
mem[4848] = 0;
mem[4849] = 0;
mem[4850] = 0;
mem[4851] = 0;
mem[4852] = 0;
mem[4853] = 0;
mem[4854] = 0;
mem[4855] = 0;
mem[4856] = 0;
mem[4857] = 0;
mem[4858] = 0;
mem[4859] = 0;

data = mem[addr];
end

endmodule